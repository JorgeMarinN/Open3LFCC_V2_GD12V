magic
tech sky130A
magscale 1 2
timestamp 1698851424
<< dnwell >>
rect -1364 -988 1364 86
<< nwell >>
rect -1370 986 -888 1318
rect -487 434 487 1368
rect 888 986 1370 1318
rect -1236 166 1236 434
rect -1444 -120 1444 166
rect -1444 -782 -1158 -120
rect 1158 -782 1444 -120
rect -1444 -1068 1444 -782
<< pwell >>
rect -1158 -782 1158 -120
<< mvnmos >>
rect -919 -502 -819 -302
rect -761 -502 -661 -302
rect -603 -502 -503 -302
rect -445 -502 -345 -302
rect -287 -502 -187 -302
rect -129 -502 -29 -302
rect 29 -502 129 -302
rect 187 -502 287 -302
rect 345 -502 445 -302
rect 503 -502 603 -302
rect 661 -502 761 -302
rect 819 -502 919 -302
rect -84 -1990 316 -1190
rect 374 -1990 774 -1190
rect 832 -1990 1232 -1190
<< mvpmos >>
rect -1112 1052 -1012 1252
rect -1112 168 -1012 368
rect -775 168 -575 268
rect -229 168 -29 1168
rect 29 168 229 1168
rect 1012 1052 1112 1252
rect 575 168 775 268
rect 1012 168 1112 368
<< mvndiff >>
rect -977 -314 -919 -302
rect -977 -490 -965 -314
rect -931 -490 -919 -314
rect -977 -502 -919 -490
rect -819 -314 -761 -302
rect -819 -490 -807 -314
rect -773 -490 -761 -314
rect -819 -502 -761 -490
rect -661 -314 -603 -302
rect -661 -490 -649 -314
rect -615 -490 -603 -314
rect -661 -502 -603 -490
rect -503 -314 -445 -302
rect -503 -490 -491 -314
rect -457 -490 -445 -314
rect -503 -502 -445 -490
rect -345 -314 -287 -302
rect -345 -490 -333 -314
rect -299 -490 -287 -314
rect -345 -502 -287 -490
rect -187 -314 -129 -302
rect -187 -490 -175 -314
rect -141 -490 -129 -314
rect -187 -502 -129 -490
rect -29 -314 29 -302
rect -29 -490 -17 -314
rect 17 -490 29 -314
rect -29 -502 29 -490
rect 129 -314 187 -302
rect 129 -490 141 -314
rect 175 -490 187 -314
rect 129 -502 187 -490
rect 287 -314 345 -302
rect 287 -490 299 -314
rect 333 -490 345 -314
rect 287 -502 345 -490
rect 445 -314 503 -302
rect 445 -490 457 -314
rect 491 -490 503 -314
rect 445 -502 503 -490
rect 603 -314 661 -302
rect 603 -490 615 -314
rect 649 -490 661 -314
rect 603 -502 661 -490
rect 761 -314 819 -302
rect 761 -490 773 -314
rect 807 -490 819 -314
rect 761 -502 819 -490
rect 919 -314 977 -302
rect 919 -490 931 -314
rect 965 -490 977 -314
rect 919 -502 977 -490
rect -142 -1202 -84 -1190
rect -142 -1978 -130 -1202
rect -96 -1978 -84 -1202
rect -142 -1990 -84 -1978
rect 316 -1202 374 -1190
rect 316 -1978 328 -1202
rect 362 -1978 374 -1202
rect 316 -1990 374 -1978
rect 774 -1202 832 -1190
rect 774 -1978 786 -1202
rect 820 -1978 832 -1202
rect 774 -1990 832 -1978
rect 1232 -1202 1290 -1190
rect 1232 -1978 1244 -1202
rect 1278 -1978 1290 -1202
rect 1232 -1990 1290 -1978
<< mvpdiff >>
rect -1170 1240 -1112 1252
rect -1170 1064 -1158 1240
rect -1124 1064 -1112 1240
rect -1170 1052 -1112 1064
rect -1012 1240 -954 1252
rect -1012 1064 -1000 1240
rect -966 1064 -954 1240
rect 954 1240 1012 1252
rect -1012 1052 -954 1064
rect -1170 356 -1112 368
rect -1170 180 -1158 356
rect -1124 180 -1112 356
rect -1170 168 -1112 180
rect -1012 356 -954 368
rect -1012 180 -1000 356
rect -966 180 -954 356
rect -1012 168 -954 180
rect -833 256 -775 268
rect -833 180 -821 256
rect -787 180 -775 256
rect -833 168 -775 180
rect -575 256 -517 268
rect -575 180 -563 256
rect -529 180 -517 256
rect -575 168 -517 180
rect -287 1156 -229 1168
rect -287 180 -275 1156
rect -241 180 -229 1156
rect -287 168 -229 180
rect -29 1156 29 1168
rect -29 180 -17 1156
rect 17 180 29 1156
rect -29 168 29 180
rect 229 1156 287 1168
rect 229 180 241 1156
rect 275 180 287 1156
rect 229 168 287 180
rect 954 1064 966 1240
rect 1000 1064 1012 1240
rect 954 1052 1012 1064
rect 1112 1240 1170 1252
rect 1112 1064 1124 1240
rect 1158 1064 1170 1240
rect 1112 1052 1170 1064
rect 954 356 1012 368
rect 517 256 575 268
rect 517 180 529 256
rect 563 180 575 256
rect 517 168 575 180
rect 775 256 833 268
rect 775 180 787 256
rect 821 180 833 256
rect 775 168 833 180
rect 954 180 966 356
rect 1000 180 1012 356
rect 954 168 1012 180
rect 1112 356 1170 368
rect 1112 180 1124 356
rect 1158 180 1170 356
rect 1112 168 1170 180
<< mvndiffc >>
rect -965 -490 -931 -314
rect -807 -490 -773 -314
rect -649 -490 -615 -314
rect -491 -490 -457 -314
rect -333 -490 -299 -314
rect -175 -490 -141 -314
rect -17 -490 17 -314
rect 141 -490 175 -314
rect 299 -490 333 -314
rect 457 -490 491 -314
rect 615 -490 649 -314
rect 773 -490 807 -314
rect 931 -490 965 -314
rect -130 -1978 -96 -1202
rect 328 -1978 362 -1202
rect 786 -1978 820 -1202
rect 1244 -1978 1278 -1202
<< mvpdiffc >>
rect -1158 1064 -1124 1240
rect -1000 1064 -966 1240
rect -1158 180 -1124 356
rect -1000 180 -966 356
rect -821 180 -787 256
rect -563 180 -529 256
rect -275 180 -241 1156
rect -17 180 17 1156
rect 241 180 275 1156
rect 966 1064 1000 1240
rect 1124 1064 1158 1240
rect 529 180 563 256
rect 787 180 821 256
rect 966 180 1000 356
rect 1124 180 1158 356
<< mvpsubdiff >>
rect -977 -168 977 -148
rect -977 -208 -947 -168
rect 947 -208 977 -168
rect -977 -228 977 -208
rect -1131 -332 -1051 -302
rect -1131 -472 -1111 -332
rect -1071 -472 -1051 -332
rect -1131 -502 -1051 -472
rect 1051 -332 1131 -302
rect 1051 -472 1071 -332
rect 1111 -472 1131 -332
rect 1051 -502 1131 -472
rect -977 -694 977 -674
rect -977 -734 -947 -694
rect 947 -734 977 -694
rect -977 -754 977 -734
rect -296 -1220 -216 -1190
rect -296 -1960 -276 -1220
rect -236 -1960 -216 -1220
rect -296 -1990 -216 -1960
rect 1364 -1220 1444 -1190
rect 1364 -1960 1384 -1220
rect 1424 -1960 1444 -1220
rect 1364 -1990 1444 -1960
rect -142 -2084 1290 -2064
rect -142 -2124 -112 -2084
rect 1260 -2124 1290 -2084
rect -142 -2144 1290 -2124
<< mvnsubdiff >>
rect -287 1282 287 1302
rect -1304 1222 -1224 1252
rect -1304 1082 -1284 1222
rect -1244 1082 -1224 1222
rect -1304 1052 -1224 1082
rect -287 1242 -257 1282
rect 257 1242 287 1282
rect -287 1222 287 1242
rect -421 1138 -341 1168
rect -421 198 -401 1138
rect -361 198 -341 1138
rect -421 168 -341 198
rect 341 1138 421 1168
rect 341 198 361 1138
rect 401 198 421 1138
rect 1224 1222 1304 1252
rect 1224 1082 1244 1222
rect 1284 1082 1304 1222
rect 1224 1052 1304 1082
rect 341 168 421 198
rect -1364 -150 -1284 -120
rect -1364 -752 -1344 -150
rect -1304 -752 -1284 -150
rect 1284 -150 1364 -120
rect -1364 -782 -1284 -752
rect 1284 -752 1304 -150
rect 1344 -752 1364 -150
rect 1284 -782 1364 -752
rect -1158 -928 1158 -908
rect -1158 -968 -1128 -928
rect 1128 -968 1158 -928
rect -1158 -988 1158 -968
<< mvpsubdiffcont >>
rect -947 -208 947 -168
rect -1111 -472 -1071 -332
rect 1071 -472 1111 -332
rect -947 -734 947 -694
rect -276 -1960 -236 -1220
rect 1384 -1960 1424 -1220
rect -112 -2124 1260 -2084
<< mvnsubdiffcont >>
rect -1284 1082 -1244 1222
rect -257 1242 257 1282
rect -401 198 -361 1138
rect 361 198 401 1138
rect 1244 1082 1284 1222
rect -1344 -752 -1304 -150
rect 1304 -752 1344 -150
rect -1128 -968 1128 -928
<< poly >>
rect -1112 1252 -1012 1278
rect 1012 1252 1112 1278
rect -229 1168 -29 1194
rect 29 1168 229 1194
rect -1112 960 -1012 1052
rect -1112 900 -1092 960
rect -1032 900 -1012 960
rect -1112 880 -1012 900
rect -1112 368 -1012 394
rect -775 268 -575 294
rect 1012 960 1112 1052
rect 1012 900 1032 960
rect 1092 900 1112 960
rect 1012 880 1112 900
rect 1012 368 1112 394
rect 575 268 775 294
rect -1112 94 -1012 168
rect -775 142 -575 168
rect -229 142 -29 168
rect 29 142 229 168
rect 575 142 775 168
rect -1112 34 -1092 94
rect -1032 34 -1012 94
rect -1112 14 -1012 34
rect -753 94 -597 142
rect -753 34 -733 94
rect -617 34 -597 94
rect -753 14 -597 34
rect -207 94 -51 142
rect -207 34 -187 94
rect -71 34 -51 94
rect -207 14 -51 34
rect 51 94 207 142
rect 51 34 71 94
rect 187 34 207 94
rect 51 14 207 34
rect 597 94 753 142
rect 597 34 617 94
rect 733 34 753 94
rect 597 14 753 34
rect 1012 94 1112 168
rect 1012 34 1032 94
rect 1092 34 1112 94
rect 1012 14 1112 34
rect -919 -302 -819 -276
rect -761 -302 -661 -276
rect -603 -302 -503 -276
rect -445 -302 -345 -276
rect -287 -302 -187 -276
rect -129 -302 -29 -276
rect 29 -302 129 -276
rect 187 -302 287 -276
rect 345 -302 445 -276
rect 503 -302 603 -276
rect 661 -302 761 -276
rect 819 -302 919 -276
rect -919 -540 -819 -502
rect -761 -540 -661 -502
rect -919 -560 -661 -540
rect -919 -620 -899 -560
rect -681 -620 -661 -560
rect -919 -640 -661 -620
rect -603 -540 -503 -502
rect -445 -540 -345 -502
rect -603 -560 -345 -540
rect -603 -620 -583 -560
rect -365 -620 -345 -560
rect -603 -640 -345 -620
rect -287 -540 -187 -502
rect -129 -540 -29 -502
rect -287 -560 -29 -540
rect -287 -620 -267 -560
rect -49 -620 -29 -560
rect -287 -640 -29 -620
rect 29 -540 129 -502
rect 187 -540 287 -502
rect 29 -560 287 -540
rect 29 -620 49 -560
rect 267 -620 287 -560
rect 29 -640 287 -620
rect 345 -540 445 -502
rect 503 -540 603 -502
rect 345 -560 603 -540
rect 345 -620 365 -560
rect 583 -620 603 -560
rect 345 -640 603 -620
rect 661 -540 761 -502
rect 819 -540 919 -502
rect 661 -560 919 -540
rect 661 -620 681 -560
rect 899 -620 919 -560
rect 661 -640 919 -620
rect -34 -1082 266 -1062
rect -34 -1142 -14 -1082
rect 246 -1142 266 -1082
rect -34 -1164 266 -1142
rect 424 -1082 724 -1062
rect 424 -1142 444 -1082
rect 704 -1142 724 -1082
rect 424 -1164 724 -1142
rect 882 -1082 1182 -1062
rect 882 -1142 902 -1082
rect 1162 -1142 1182 -1082
rect 882 -1164 1182 -1142
rect -84 -1190 316 -1164
rect 374 -1190 774 -1164
rect 832 -1190 1232 -1164
rect -84 -2016 316 -1990
rect 374 -2016 774 -1990
rect 832 -2016 1232 -1990
<< polycont >>
rect -1092 900 -1032 960
rect 1032 900 1092 960
rect -1092 34 -1032 94
rect -733 34 -617 94
rect -187 34 -71 94
rect 71 34 187 94
rect 617 34 733 94
rect 1032 34 1092 94
rect -899 -620 -681 -560
rect -583 -620 -365 -560
rect -267 -620 -49 -560
rect 49 -620 267 -560
rect 365 -620 583 -560
rect 681 -620 899 -560
rect -14 -1142 246 -1082
rect 444 -1142 704 -1082
rect 902 -1142 1162 -1082
<< locali >>
rect -287 1282 287 1302
rect -1304 1222 -1224 1252
rect -1304 1082 -1284 1222
rect -1244 1082 -1224 1222
rect -1304 1052 -1224 1082
rect -1158 1240 -1124 1256
rect -1158 1048 -1124 1064
rect -1000 1240 -966 1256
rect -287 1242 -257 1282
rect 257 1242 287 1282
rect -287 1222 287 1242
rect 966 1240 1000 1256
rect -1000 1048 -966 1064
rect -421 1138 -341 1168
rect -1112 960 -954 980
rect -1112 900 -1092 960
rect -974 900 -954 960
rect -1112 880 -954 900
rect -1158 356 -1124 372
rect -1158 164 -1124 180
rect -1000 356 -966 372
rect -1000 164 -966 180
rect -821 256 -787 272
rect -821 164 -787 180
rect -563 256 -529 272
rect -563 164 -529 180
rect -421 198 -401 1138
rect -361 198 -341 1138
rect -421 168 -341 198
rect -275 1156 -241 1172
rect -275 164 -241 180
rect -17 1156 17 1172
rect -17 164 17 180
rect 241 1156 275 1172
rect 241 164 275 180
rect 341 1138 421 1168
rect 341 198 361 1138
rect 401 198 421 1138
rect 966 1048 1000 1064
rect 1124 1240 1158 1256
rect 1124 1048 1158 1064
rect 1224 1222 1304 1252
rect 1224 1082 1244 1222
rect 1284 1082 1304 1222
rect 1224 1052 1304 1082
rect 954 960 1112 980
rect 954 900 974 960
rect 1092 900 1112 960
rect 954 880 1112 900
rect 966 356 1000 372
rect 341 168 421 198
rect 529 256 563 272
rect 529 164 563 180
rect 787 256 821 272
rect 787 164 821 180
rect 966 164 1000 180
rect 1124 356 1158 372
rect 1124 164 1158 180
rect -1112 94 -1012 114
rect -1112 34 -1092 94
rect -1032 34 -1012 94
rect -1112 14 -1012 34
rect -753 94 -597 114
rect -753 34 -733 94
rect -617 34 -597 94
rect -753 -34 -597 34
rect -753 -94 -733 -34
rect -617 -94 -597 -34
rect -753 -114 -597 -94
rect -207 94 -51 114
rect -207 34 -187 94
rect -71 34 -51 94
rect -207 -34 -51 34
rect 51 94 207 114
rect 51 34 71 94
rect 187 34 207 94
rect 51 14 207 34
rect 597 94 753 114
rect 597 34 617 94
rect 733 34 753 94
rect 597 14 753 34
rect 1012 94 1112 114
rect 1012 34 1032 94
rect 1092 34 1112 94
rect -207 -94 -187 -34
rect -71 -94 -51 -34
rect -207 -114 -51 -94
rect 1012 -34 1112 34
rect 1012 -94 1032 -34
rect 1092 -94 1112 -34
rect 1012 -114 1112 -94
rect -1364 -150 -1284 -120
rect -1364 -752 -1344 -150
rect -1304 -752 -1284 -150
rect -1131 -168 1131 -148
rect -1131 -208 -947 -168
rect 947 -208 1131 -168
rect -1131 -228 1131 -208
rect -1131 -332 -1051 -228
rect -1131 -472 -1111 -332
rect -1071 -472 -1051 -332
rect -1131 -502 -1051 -472
rect -965 -314 -931 -298
rect -965 -506 -931 -490
rect -807 -314 -773 -298
rect -807 -506 -773 -490
rect -649 -314 -615 -298
rect -649 -506 -615 -490
rect -491 -314 -457 -298
rect -491 -506 -457 -490
rect -333 -314 -299 -298
rect -333 -506 -299 -490
rect -175 -314 -141 -298
rect -175 -506 -141 -490
rect -17 -314 17 -298
rect -17 -506 17 -490
rect 141 -314 175 -298
rect 141 -506 175 -490
rect 299 -314 333 -298
rect 299 -506 333 -490
rect 457 -314 491 -298
rect 457 -506 491 -490
rect 615 -314 649 -298
rect 615 -506 649 -490
rect 773 -314 807 -298
rect 773 -506 807 -490
rect 931 -314 965 -298
rect 931 -506 965 -490
rect 1051 -332 1131 -228
rect 1051 -472 1071 -332
rect 1111 -472 1131 -332
rect 1051 -502 1131 -472
rect 1284 -150 1364 -120
rect -919 -560 -661 -540
rect -919 -620 -899 -560
rect -681 -620 -661 -560
rect -919 -640 -661 -620
rect -603 -560 -345 -540
rect -603 -620 -583 -560
rect -365 -620 -345 -560
rect -603 -640 -345 -620
rect -287 -560 -29 -540
rect -287 -620 -267 -560
rect -49 -620 -29 -560
rect -287 -640 -29 -620
rect 29 -560 287 -540
rect 29 -620 49 -560
rect 267 -620 287 -560
rect 29 -640 287 -620
rect 345 -560 603 -540
rect 345 -620 365 -560
rect 583 -620 603 -560
rect 345 -640 603 -620
rect 661 -560 919 -540
rect 661 -620 681 -560
rect 899 -620 919 -560
rect 661 -640 919 -620
rect -1364 -782 -1284 -752
rect -977 -694 977 -674
rect -977 -734 -947 -694
rect 947 -734 977 -694
rect -977 -754 977 -734
rect 1284 -752 1304 -150
rect 1344 -752 1364 -150
rect 1284 -782 1364 -752
rect -1158 -928 1158 -908
rect -1158 -968 -1128 -928
rect 1128 -968 1158 -928
rect -1158 -988 1158 -968
rect -34 -1082 266 -1062
rect -34 -1142 -14 -1082
rect 246 -1142 266 -1082
rect -34 -1162 266 -1142
rect 424 -1082 724 -1062
rect 424 -1142 444 -1082
rect 704 -1142 724 -1082
rect 424 -1162 724 -1142
rect 882 -1082 1182 -1062
rect 882 -1142 902 -1082
rect 1162 -1142 1182 -1082
rect 882 -1162 1182 -1142
rect -296 -1220 -216 -1190
rect -296 -1960 -276 -1220
rect -236 -1960 -216 -1220
rect -296 -1990 -216 -1960
rect -130 -1202 -96 -1186
rect -130 -1994 -96 -1978
rect 328 -1202 362 -1186
rect 328 -1994 362 -1978
rect 786 -1202 820 -1186
rect 786 -1994 820 -1978
rect 1244 -1202 1278 -1186
rect 1244 -1994 1278 -1978
rect 1364 -1220 1444 -1190
rect 1364 -1960 1384 -1220
rect 1424 -1960 1444 -1220
rect 1364 -1990 1444 -1960
rect -142 -2084 1290 -2064
rect -142 -2124 -112 -2084
rect 1260 -2124 1290 -2084
rect -142 -2144 1290 -2124
<< viali >>
rect -1284 1082 -1244 1222
rect -1158 1064 -1124 1240
rect -1000 1064 -966 1240
rect -257 1242 257 1282
rect -1034 900 -1032 960
rect -1032 900 -974 960
rect -1158 180 -1124 356
rect -1000 180 -966 356
rect -821 180 -787 256
rect -563 180 -529 256
rect -401 198 -361 1138
rect -275 180 -241 1156
rect -17 180 17 1156
rect 241 180 275 1156
rect 361 198 401 1138
rect 966 1064 1000 1240
rect 1124 1064 1158 1240
rect 1244 1082 1284 1222
rect 974 900 1032 960
rect 1032 900 1034 960
rect 529 180 563 256
rect 787 180 821 256
rect 966 180 1000 356
rect 1124 180 1158 356
rect -1092 34 -1032 94
rect -733 -94 -617 -34
rect 71 34 187 94
rect 617 34 733 94
rect -187 -94 -71 -34
rect 1032 -94 1092 -34
rect -1344 -752 -1304 -150
rect -1111 -472 -1071 -332
rect -965 -490 -931 -314
rect -807 -490 -773 -314
rect -649 -490 -615 -314
rect -491 -490 -457 -314
rect -333 -490 -299 -314
rect -175 -490 -141 -314
rect -17 -490 17 -314
rect 141 -490 175 -314
rect 299 -490 333 -314
rect 457 -490 491 -314
rect 615 -490 649 -314
rect 773 -490 807 -314
rect 931 -490 965 -314
rect 1071 -472 1111 -332
rect -877 -620 -703 -560
rect -561 -620 -387 -560
rect -245 -620 -71 -560
rect 71 -620 245 -560
rect 387 -620 561 -560
rect 703 -620 877 -560
rect -947 -734 947 -694
rect 1304 -752 1344 -150
rect -1128 -968 670 -928
rect 930 -968 1128 -928
rect -14 -1142 246 -1082
rect 444 -1142 704 -1082
rect 902 -1142 1162 -1082
rect -276 -1960 -236 -1220
rect -130 -1978 -96 -1202
rect 328 -1978 362 -1202
rect 786 -1978 820 -1202
rect 1244 -1978 1278 -1202
rect 1384 -1960 1424 -1220
rect -112 -2124 1260 -2084
<< metal1 >>
rect -441 1282 441 1422
rect -1304 1240 -1118 1252
rect -1304 1222 -1158 1240
rect -1304 1082 -1284 1222
rect -1244 1082 -1158 1222
rect -1304 1064 -1158 1082
rect -1124 1064 -1118 1240
rect -1304 1052 -1118 1064
rect -1384 528 -1284 548
rect -1384 468 -1364 528
rect -1304 468 -1284 528
rect -1384 -150 -1284 468
rect -1164 356 -1118 1052
rect -1006 1240 -960 1252
rect -1006 1064 -1000 1240
rect -966 1064 -960 1240
rect -1006 980 -960 1064
rect -441 1242 -257 1282
rect 257 1242 441 1282
rect -441 1222 441 1242
rect -441 1138 -341 1222
rect -1090 960 -469 980
rect -1090 900 -1034 960
rect -974 900 -469 960
rect -1090 880 -469 900
rect -1164 180 -1158 356
rect -1124 180 -1118 356
rect -1164 168 -1118 180
rect -1006 528 -781 548
rect -1006 468 -986 528
rect -801 468 -781 528
rect -1006 356 -781 468
rect -1006 180 -1000 356
rect -966 256 -781 356
rect -966 180 -821 256
rect -787 180 -781 256
rect -1006 168 -781 180
rect -569 256 -469 880
rect -569 180 -563 256
rect -529 180 -469 256
rect -1112 94 -1012 114
rect -1112 34 -1092 94
rect -1032 34 -1012 94
rect -1112 14 -1012 34
rect -569 -14 -469 180
rect -441 528 -401 1138
rect -441 468 -421 528
rect -441 198 -401 468
rect -361 198 -341 1138
rect -441 168 -341 198
rect -281 1156 -235 1168
rect -281 180 -275 1156
rect -241 180 -235 1156
rect -281 114 -235 180
rect -23 1156 23 1222
rect -23 180 -17 1156
rect 17 180 23 1156
rect -23 168 23 180
rect 235 1156 281 1168
rect 235 180 241 1156
rect 275 180 281 1156
rect -308 94 -208 114
rect -308 34 -288 94
rect -228 34 -208 94
rect -308 14 -208 34
rect 51 94 207 114
rect 51 34 71 94
rect 187 34 207 94
rect 51 14 207 34
rect -840 -34 -451 -14
rect -840 -94 -820 -34
rect -760 -94 -733 -34
rect -617 -94 -549 -34
rect -489 -94 -451 -34
rect -840 -114 -451 -94
rect -207 -34 -51 -14
rect -207 -94 -187 -34
rect -71 -94 -51 -34
rect -207 -114 -51 -94
rect -1384 -752 -1344 -150
rect -1304 -752 -1284 -150
rect -1384 -908 -1284 -752
rect -1131 -314 -925 -302
rect -1131 -332 -965 -314
rect -1131 -472 -1111 -332
rect -1071 -472 -965 -332
rect -1131 -490 -965 -472
rect -931 -490 -925 -314
rect -1131 -674 -925 -490
rect -813 -314 -767 -114
rect -813 -490 -807 -314
rect -773 -490 -767 -314
rect -813 -502 -767 -490
rect -655 -314 -609 -302
rect -655 -490 -649 -314
rect -615 -490 -609 -314
rect -897 -560 -683 -540
rect -897 -620 -877 -560
rect -703 -620 -683 -560
rect -897 -640 -683 -620
rect -655 -674 -609 -490
rect -497 -314 -451 -114
rect -497 -490 -491 -314
rect -457 -490 -451 -314
rect -497 -502 -451 -490
rect -339 -314 -293 -302
rect -339 -490 -333 -314
rect -299 -490 -293 -314
rect -581 -560 -367 -540
rect -581 -620 -561 -560
rect -387 -620 -367 -560
rect -581 -640 -367 -620
rect -339 -674 -293 -490
rect -181 -314 -135 -114
rect -181 -490 -175 -314
rect -141 -490 -135 -314
rect -181 -502 -135 -490
rect -23 -314 23 -302
rect -23 -490 -17 -314
rect 17 -490 23 -314
rect -265 -560 -51 -540
rect -265 -620 -245 -560
rect -71 -620 -51 -560
rect -265 -640 -51 -620
rect -23 -674 23 -490
rect 135 -314 181 14
rect 235 -14 281 180
rect 341 1138 441 1222
rect 341 198 361 1138
rect 401 528 441 1138
rect 960 1240 1006 1252
rect 960 1064 966 1240
rect 1000 1064 1006 1240
rect 960 980 1006 1064
rect 1118 1240 1304 1252
rect 1118 1064 1124 1240
rect 1158 1222 1304 1240
rect 1158 1082 1244 1222
rect 1284 1082 1304 1222
rect 1158 1064 1304 1082
rect 1118 1052 1304 1064
rect 421 468 441 528
rect 401 198 441 468
rect 341 168 441 198
rect 469 960 1090 980
rect 469 900 974 960
rect 1034 900 1090 960
rect 469 880 1090 900
rect 469 256 569 880
rect 469 180 529 256
rect 563 180 569 256
rect 469 114 569 180
rect 781 528 1006 548
rect 781 468 801 528
rect 986 468 1006 528
rect 781 356 1006 468
rect 781 256 966 356
rect 781 180 787 256
rect 821 180 966 256
rect 1000 180 1006 356
rect 781 168 1006 180
rect 1118 356 1164 1052
rect 1118 180 1124 356
rect 1158 180 1164 356
rect 1118 168 1164 180
rect 1284 528 1384 548
rect 1284 468 1304 528
rect 1364 468 1384 528
rect 451 94 840 114
rect 451 34 489 94
rect 549 34 617 94
rect 733 34 760 94
rect 820 34 840 94
rect 451 14 840 34
rect 228 -34 328 -14
rect 228 -94 248 -34
rect 308 -94 328 -34
rect 228 -114 328 -94
rect 135 -490 141 -314
rect 175 -490 181 -314
rect 135 -502 181 -490
rect 293 -314 339 -302
rect 293 -490 299 -314
rect 333 -490 339 -314
rect 51 -560 265 -540
rect 51 -620 71 -560
rect 245 -620 265 -560
rect 51 -640 265 -620
rect 293 -674 339 -490
rect 451 -314 497 14
rect 451 -490 457 -314
rect 491 -490 497 -314
rect 451 -502 497 -490
rect 609 -314 655 -302
rect 609 -490 615 -314
rect 649 -490 655 -314
rect 367 -560 581 -540
rect 367 -620 387 -560
rect 561 -620 581 -560
rect 367 -640 581 -620
rect 609 -674 655 -490
rect 767 -314 813 14
rect 1012 -34 1112 -14
rect 1012 -94 1032 -34
rect 1092 -94 1112 -34
rect 1012 -114 1112 -94
rect 1284 -150 1384 468
rect 767 -490 773 -314
rect 807 -490 813 -314
rect 767 -502 813 -490
rect 925 -314 1131 -302
rect 925 -490 931 -314
rect 965 -332 1131 -314
rect 965 -472 1071 -332
rect 1111 -472 1131 -332
rect 965 -490 1131 -472
rect 683 -560 897 -540
rect 683 -620 703 -560
rect 877 -620 897 -560
rect 683 -640 897 -620
rect 925 -674 1131 -490
rect -1131 -694 1131 -674
rect -1131 -734 -947 -694
rect 947 -734 1131 -694
rect -1131 -774 1131 -734
rect 1284 -752 1304 -150
rect 1344 -752 1384 -150
rect -1384 -928 700 -908
rect -1384 -968 -1128 -928
rect 670 -968 700 -928
rect -1384 -1008 700 -968
rect -136 -1082 266 -1062
rect -136 -1142 -14 -1082
rect 246 -1142 266 -1082
rect -136 -1162 266 -1142
rect 424 -1082 724 -1062
rect 424 -1142 444 -1082
rect 704 -1142 724 -1082
rect 424 -1162 724 -1142
rect 753 -1162 853 -774
rect 1284 -908 1384 -752
rect 900 -928 1384 -908
rect 900 -968 930 -928
rect 1128 -968 1384 -928
rect 900 -1008 1384 -968
rect 882 -1082 1182 -1062
rect 882 -1142 902 -1082
rect 1162 -1142 1182 -1082
rect 882 -1162 1182 -1142
rect -296 -1220 -216 -1190
rect -296 -1960 -276 -1220
rect -236 -1960 -216 -1220
rect -296 -2064 -216 -1960
rect -136 -1202 -90 -1162
rect -136 -1978 -130 -1202
rect -96 -1978 -90 -1202
rect -136 -1990 -90 -1978
rect 322 -1202 368 -1190
rect 322 -1978 328 -1202
rect 362 -1978 368 -1202
rect 322 -2064 368 -1978
rect 780 -1202 826 -1162
rect 780 -1978 786 -1202
rect 820 -1978 826 -1202
rect 780 -1990 826 -1978
rect 1238 -1202 1444 -1190
rect 1238 -1978 1244 -1202
rect 1278 -1220 1444 -1202
rect 1278 -1960 1384 -1220
rect 1424 -1960 1444 -1220
rect 1278 -1978 1444 -1960
rect 1238 -1990 1444 -1978
rect 1284 -2064 1444 -1990
rect -296 -2084 1444 -2064
rect -296 -2124 -112 -2084
rect 1260 -2124 1444 -2084
rect -296 -2264 1444 -2124
<< via1 >>
rect -1364 468 -1304 528
rect -986 468 -801 528
rect -1092 34 -1032 94
rect -421 468 -401 528
rect -401 468 -361 528
rect -288 34 -228 94
rect 71 34 187 94
rect -820 -94 -760 -34
rect -733 -94 -617 -34
rect -549 -94 -489 -34
rect -187 -94 -71 -34
rect -877 -620 -703 -560
rect -561 -620 -387 -560
rect -245 -620 -71 -560
rect 361 468 401 528
rect 401 468 421 528
rect 801 468 986 528
rect 1304 468 1364 528
rect 489 34 549 94
rect 617 34 733 94
rect 760 34 820 94
rect 248 -94 308 -34
rect 71 -620 245 -560
rect 387 -620 561 -560
rect 1032 -94 1092 -34
rect 703 -620 877 -560
rect -14 -1142 246 -1082
rect 444 -1142 704 -1082
rect 902 -1142 1162 -1082
<< metal2 >>
rect -1384 528 -341 548
rect -1384 468 -1364 528
rect -1304 468 -986 528
rect -801 468 -421 528
rect -361 468 -341 528
rect -1384 448 -341 468
rect 341 528 1384 548
rect 341 468 361 528
rect 421 468 801 528
rect 986 468 1304 528
rect 1364 468 1384 528
rect 341 448 1384 468
rect -1154 94 1444 114
rect -1154 34 -1092 94
rect -1032 34 -288 94
rect -228 34 71 94
rect 187 34 489 94
rect 549 34 617 94
rect 733 34 760 94
rect 820 34 1444 94
rect -1154 14 1444 34
rect -1154 -34 1444 -14
rect -1154 -94 -820 -34
rect -760 -94 -733 -34
rect -617 -94 -549 -34
rect -489 -94 -187 -34
rect -71 -94 248 -34
rect 308 -94 1032 -34
rect 1092 -94 1444 -34
rect -1154 -114 1444 -94
rect -977 -560 -29 -540
rect -977 -620 -877 -560
rect -703 -620 -561 -560
rect -387 -620 -245 -560
rect -71 -620 -29 -560
rect -977 -640 -29 -620
rect 29 -560 977 -540
rect 29 -620 71 -560
rect 245 -620 387 -560
rect 561 -620 703 -560
rect 877 -620 977 -560
rect 29 -640 977 -620
rect -742 -1082 1210 -1062
rect -742 -1142 -14 -1082
rect 246 -1142 444 -1082
rect 704 -1142 902 -1082
rect 1162 -1142 1210 -1082
rect -742 -1162 1210 -1142
<< labels >>
rlabel metal1 -441 1322 -341 1422 1 VDD
rlabel metal2 1344 14 1444 114 3 RESET
rlabel metal2 1344 -114 1444 -14 3 SET
rlabel metal2 -977 -640 -29 -540 7 VRE
rlabel metal2 29 -640 977 -540 3 VFE
rlabel metal2 -742 -1162 -642 -1062 7 Iref
rlabel metal1 -296 -2264 -196 -2164 5 GND
<< end >>
