magic
tech sky130A
magscale 1 2
timestamp 1699989067
<< locali >>
rect 111768 -16596 113018 -16551
rect 111768 -16898 111878 -16596
rect 112876 -16898 113018 -16596
rect 111768 -16972 113018 -16898
<< viali >>
rect 111878 -16898 112876 -16596
<< metal1 >>
rect 6000 -620 6320 -600
rect 6000 -4080 6020 -620
rect 6000 -4200 6320 -4080
rect 15008 -620 15400 -600
rect 15008 -6420 15020 -620
rect 15380 -6420 15400 -620
rect 15008 -6600 15400 -6420
rect 4000 -6820 9600 -6800
rect 4000 -7180 9220 -6820
rect 9580 -7180 9600 -6820
rect 4000 -7200 9600 -7180
rect 6000 -10020 112000 -10000
rect 6000 -10380 6020 -10020
rect 6380 -10380 112000 -10020
rect 6000 -10400 112000 -10380
rect 112220 -12800 112320 -12780
rect 112220 -13200 112240 -12800
rect 112300 -13200 112320 -12800
rect 112220 -13220 112320 -13200
rect 110839 -14667 111871 -14525
rect 110839 -15736 110913 -14667
rect 111200 -15736 111871 -14667
rect 110839 -15852 111871 -15736
rect 111784 -16596 112953 -16547
rect 111784 -16898 111878 -16596
rect 112876 -16898 112953 -16596
rect 111784 -16962 112953 -16898
rect 9200 -44820 112000 -44800
rect 9200 -45180 9220 -44820
rect 9580 -45180 112000 -44820
rect 9200 -45200 112000 -45180
rect 15000 -45420 112400 -45400
rect 15000 -46380 15020 -45420
rect 15380 -46380 112240 -45420
rect 112300 -46380 112400 -45420
rect 15000 -46400 112400 -46380
<< via1 >>
rect 6020 -4080 6320 -620
rect 9400 -6000 9454 -5500
rect 15020 -6420 15380 -620
rect 9220 -7180 9580 -6820
rect 6020 -10380 6380 -10020
rect 112240 -13200 112300 -12800
rect 110913 -15736 111200 -14667
rect 112066 -16827 112642 -16647
rect 9220 -45180 9580 -44820
rect 15020 -46380 15380 -45420
rect 112240 -46380 112300 -45420
<< metal2 >>
rect 58000 56000 66000 60000
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 6000 580 6400 600
rect 6000 20 6020 580
rect 6380 20 6400 580
rect 6000 -620 6400 20
rect 6000 -4080 6020 -620
rect 6320 -4080 6400 -620
rect 10434 -800 10754 5440
rect 58000 2000 66000 6000
rect 15000 -620 15400 -600
rect 6000 -10020 6400 -4080
rect 9384 -6000 9400 -5500
rect 9454 -6000 9470 -5500
rect 9384 -6800 9470 -6000
rect 15000 -6420 15020 -620
rect 15380 -6420 15400 -620
rect 6000 -10380 6020 -10020
rect 6380 -10380 6400 -10020
rect 6000 -10400 6400 -10380
rect 9200 -6820 9600 -6800
rect 9200 -7180 9220 -6820
rect 9580 -7180 9600 -6820
rect 9200 -44820 9600 -7180
rect 9200 -45180 9220 -44820
rect 9580 -45180 9600 -44820
rect 9200 -45200 9600 -45180
rect 15000 -45420 15400 -6420
rect 112220 -12800 112320 -12780
rect 112220 -13200 112240 -12800
rect 112300 -13200 112320 -12800
rect 110839 -14667 111272 -14528
rect 110839 -15736 110913 -14667
rect 111200 -15736 111272 -14667
rect 110839 -15852 111272 -15736
rect 112220 -16580 112320 -13200
rect 111985 -16647 112726 -16580
rect 111985 -16827 112066 -16647
rect 112642 -16827 112726 -16647
rect 111985 -16895 112726 -16827
rect 15000 -46380 15020 -45420
rect 15380 -46380 15400 -45420
rect 15000 -46400 15400 -46380
rect 112220 -45420 112320 -16895
rect 112220 -46380 112240 -45420
rect 112300 -46380 112320 -45420
rect 112220 -46400 112320 -46380
<< via2 >>
rect 116000 54000 120000 58000
rect 10474 5440 10714 6360
rect 6020 20 6380 580
rect 110913 -15736 111200 -14667
<< metal3 >>
rect 6000 580 6400 12000
rect 6000 20 6020 580
rect 6380 20 6400 580
rect 6000 0 6400 20
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 10434 -800 10754 5440
rect 22000 1560 108000 1600
rect 22000 440 22040 1560
rect 107960 440 108000 1560
rect 22000 0 108000 440
rect 110000 -2040 111400 -2000
rect 110000 -43960 110040 -2040
rect 111360 -43960 111400 -2040
rect 110000 -44000 111400 -43960
<< via3 >>
rect 116000 54000 120000 58000
rect 10474 5440 10714 6360
rect 22040 440 107960 1560
rect 110040 -14667 111360 -2040
rect 110040 -15736 110913 -14667
rect 110913 -15736 111200 -14667
rect 111200 -15736 111360 -14667
rect 110040 -43960 111360 -15736
<< metal4 >>
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 10434 -800 10754 5440
rect 22000 1560 108000 2000
rect 22000 440 22040 1560
rect 107960 440 108000 1560
rect 22000 400 108000 440
rect 109320 -2040 111400 -2000
rect 109320 -43960 110040 -2040
rect 111360 -43960 111400 -2040
rect 109320 -44000 111400 -43960
<< via4 >>
rect 116000 54000 120000 58000
rect 10474 5440 10714 6360
rect 22040 440 107960 1560
<< metal5 >>
rect 2000 56000 6000 60000
rect 116000 58000 120000 60000
rect 60000 46000 64000 50000
rect 10434 6360 10754 6400
rect 10434 5440 10474 6360
rect 10714 5440 10754 6360
rect 10434 -800 10754 5440
rect 22000 1560 108000 1600
rect 22000 440 22040 1560
rect 107960 440 108000 1560
rect 22000 0 108000 440
use driver_bootstrap  driver_bootstrap_0
timestamp 1699974556
transform 0 1 113012 1 0 -8631
box -4589 -1612 7801 2600
use level_shifter  level_shifter_0
timestamp 1666543010
transform 0 1 6200 1 0 -6600
box 0 0 6050 8936
use mimcap_210x420  mimcap_210x420_0
timestamp 1698868607
transform 1 0 20000 0 1 -44660
box 0 0 89320 44660
use power_stage_3  power_stage_3_0
timestamp 1699898483
transform 0 1 0 1 0 0
box 0 0 61200 123200
use pw2nd_diode_12u7_12u7  pw2nd_diode_12u7_12u7_0
timestamp 1699972156
transform 1 0 111653 0 1 -16547
box -53 -53 2763 2763
<< labels >>
rlabel metal5 2000 56000 6000 60000 1 VSS
rlabel metal5 116000 56000 120000 60000 1 VDD
rlabel metal5 60000 46000 64000 50000 1 Vout
<< end >>
