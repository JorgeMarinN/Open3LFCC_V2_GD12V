magic
tech sky130A
timestamp 1698510666
<< nwell >>
rect 203 558 1836 1325
rect -87 112 1836 558
rect 203 107 1836 112
<< mvnmos >>
rect 29 -309 79 -9
rect 108 -309 158 -9
rect 323 -413 373 -13
rect 402 -413 452 -13
rect 481 -413 531 -13
rect 560 -413 610 -13
rect 639 -413 689 -13
rect 718 -413 768 -13
rect 797 -413 847 -13
rect 876 -413 926 -13
rect 955 -413 1005 -13
rect 1034 -413 1084 -13
rect 1113 -413 1163 -13
rect 1192 -413 1242 -13
rect 1271 -413 1321 -13
rect 1350 -413 1400 -13
rect 1429 -413 1479 -13
rect 1508 -413 1558 -13
rect 1587 -413 1637 -13
rect 1666 -413 1716 -13
<< mvpmos >>
rect 29 145 79 445
rect 108 145 158 445
rect 323 140 373 1224
rect 402 140 452 1224
rect 481 140 531 1224
rect 560 140 610 1224
rect 639 140 689 1224
rect 718 140 768 1224
rect 797 140 847 1224
rect 876 140 926 1224
rect 955 140 1005 1224
rect 1034 140 1084 1224
rect 1113 140 1163 1224
rect 1192 140 1242 1224
rect 1271 140 1321 1224
rect 1350 140 1400 1224
rect 1429 140 1479 1224
rect 1508 140 1558 1224
rect 1587 140 1637 1224
rect 1666 140 1716 1224
<< mvndiff >>
rect 0 -15 29 -9
rect 0 -303 6 -15
rect 23 -303 29 -15
rect 0 -309 29 -303
rect 79 -15 108 -9
rect 79 -303 85 -15
rect 102 -303 108 -15
rect 79 -309 108 -303
rect 158 -15 187 -9
rect 158 -303 164 -15
rect 181 -303 187 -15
rect 158 -309 187 -303
rect 294 -19 323 -13
rect 294 -407 300 -19
rect 317 -407 323 -19
rect 294 -413 323 -407
rect 373 -19 402 -13
rect 373 -407 379 -19
rect 396 -407 402 -19
rect 373 -413 402 -407
rect 452 -19 481 -13
rect 452 -407 458 -19
rect 475 -407 481 -19
rect 452 -413 481 -407
rect 531 -19 560 -13
rect 531 -407 537 -19
rect 554 -407 560 -19
rect 531 -413 560 -407
rect 610 -19 639 -13
rect 610 -407 616 -19
rect 633 -407 639 -19
rect 610 -413 639 -407
rect 689 -19 718 -13
rect 689 -407 695 -19
rect 712 -407 718 -19
rect 689 -413 718 -407
rect 768 -19 797 -13
rect 768 -407 774 -19
rect 791 -407 797 -19
rect 768 -413 797 -407
rect 847 -19 876 -13
rect 847 -407 853 -19
rect 870 -407 876 -19
rect 847 -413 876 -407
rect 926 -19 955 -13
rect 926 -407 932 -19
rect 949 -407 955 -19
rect 926 -413 955 -407
rect 1005 -19 1034 -13
rect 1005 -407 1011 -19
rect 1028 -407 1034 -19
rect 1005 -413 1034 -407
rect 1084 -19 1113 -13
rect 1084 -407 1090 -19
rect 1107 -407 1113 -19
rect 1084 -413 1113 -407
rect 1163 -19 1192 -13
rect 1163 -407 1169 -19
rect 1186 -407 1192 -19
rect 1163 -413 1192 -407
rect 1242 -19 1271 -13
rect 1242 -407 1248 -19
rect 1265 -407 1271 -19
rect 1242 -413 1271 -407
rect 1321 -19 1350 -13
rect 1321 -407 1327 -19
rect 1344 -407 1350 -19
rect 1321 -413 1350 -407
rect 1400 -19 1429 -13
rect 1400 -407 1406 -19
rect 1423 -407 1429 -19
rect 1400 -413 1429 -407
rect 1479 -19 1508 -13
rect 1479 -407 1485 -19
rect 1502 -407 1508 -19
rect 1479 -413 1508 -407
rect 1558 -19 1587 -13
rect 1558 -407 1564 -19
rect 1581 -407 1587 -19
rect 1558 -413 1587 -407
rect 1637 -19 1666 -13
rect 1637 -407 1643 -19
rect 1660 -407 1666 -19
rect 1637 -413 1666 -407
rect 1716 -19 1745 -13
rect 1716 -407 1722 -19
rect 1739 -407 1745 -19
rect 1716 -413 1745 -407
<< mvpdiff >>
rect 0 439 29 445
rect 0 151 6 439
rect 23 151 29 439
rect 0 145 29 151
rect 79 439 108 445
rect 79 151 85 439
rect 102 151 108 439
rect 79 145 108 151
rect 158 439 187 445
rect 158 151 164 439
rect 181 151 187 439
rect 158 145 187 151
rect 294 1218 323 1224
rect 294 146 300 1218
rect 317 146 323 1218
rect 294 140 323 146
rect 373 1218 402 1224
rect 373 146 379 1218
rect 396 146 402 1218
rect 373 140 402 146
rect 452 1218 481 1224
rect 452 146 458 1218
rect 475 146 481 1218
rect 452 140 481 146
rect 531 1218 560 1224
rect 531 146 537 1218
rect 554 146 560 1218
rect 531 140 560 146
rect 610 1218 639 1224
rect 610 146 616 1218
rect 633 146 639 1218
rect 610 140 639 146
rect 689 1218 718 1224
rect 689 146 695 1218
rect 712 146 718 1218
rect 689 140 718 146
rect 768 1218 797 1224
rect 768 146 774 1218
rect 791 146 797 1218
rect 768 140 797 146
rect 847 1218 876 1224
rect 847 146 853 1218
rect 870 146 876 1218
rect 847 140 876 146
rect 926 1218 955 1224
rect 926 146 932 1218
rect 949 146 955 1218
rect 926 140 955 146
rect 1005 1218 1034 1224
rect 1005 146 1011 1218
rect 1028 146 1034 1218
rect 1005 140 1034 146
rect 1084 1218 1113 1224
rect 1084 146 1090 1218
rect 1107 146 1113 1218
rect 1084 140 1113 146
rect 1163 1218 1192 1224
rect 1163 146 1169 1218
rect 1186 146 1192 1218
rect 1163 140 1192 146
rect 1242 1218 1271 1224
rect 1242 146 1248 1218
rect 1265 146 1271 1218
rect 1242 140 1271 146
rect 1321 1218 1350 1224
rect 1321 146 1327 1218
rect 1344 146 1350 1218
rect 1321 140 1350 146
rect 1400 1218 1429 1224
rect 1400 146 1406 1218
rect 1423 146 1429 1218
rect 1400 140 1429 146
rect 1479 1218 1508 1224
rect 1479 146 1485 1218
rect 1502 146 1508 1218
rect 1479 140 1508 146
rect 1558 1218 1587 1224
rect 1558 146 1564 1218
rect 1581 146 1587 1218
rect 1558 140 1587 146
rect 1637 1218 1666 1224
rect 1637 146 1643 1218
rect 1660 146 1666 1218
rect 1637 140 1666 146
rect 1716 1218 1745 1224
rect 1716 146 1722 1218
rect 1739 146 1745 1218
rect 1716 140 1745 146
<< mvndiffc >>
rect 6 -303 23 -15
rect 85 -303 102 -15
rect 164 -303 181 -15
rect 300 -407 317 -19
rect 379 -407 396 -19
rect 458 -407 475 -19
rect 537 -407 554 -19
rect 616 -407 633 -19
rect 695 -407 712 -19
rect 774 -407 791 -19
rect 853 -407 870 -19
rect 932 -407 949 -19
rect 1011 -407 1028 -19
rect 1090 -407 1107 -19
rect 1169 -407 1186 -19
rect 1248 -407 1265 -19
rect 1327 -407 1344 -19
rect 1406 -407 1423 -19
rect 1485 -407 1502 -19
rect 1564 -407 1581 -19
rect 1643 -407 1660 -19
rect 1722 -407 1739 -19
<< mvpdiffc >>
rect 6 151 23 439
rect 85 151 102 439
rect 164 151 181 439
rect 300 146 317 1218
rect 379 146 396 1218
rect 458 146 475 1218
rect 537 146 554 1218
rect 616 146 633 1218
rect 695 146 712 1218
rect 774 146 791 1218
rect 853 146 870 1218
rect 932 146 949 1218
rect 1011 146 1028 1218
rect 1090 146 1107 1218
rect 1169 146 1186 1218
rect 1248 146 1265 1218
rect 1327 146 1344 1218
rect 1406 146 1423 1218
rect 1485 146 1502 1218
rect 1564 146 1581 1218
rect 1643 146 1660 1218
rect 1722 146 1739 1218
<< mvpsubdiff >>
rect -54 -29 -37 -9
rect -54 -309 -37 -289
rect 236 -30 257 -13
rect 236 -413 257 -383
rect 1782 -30 1803 -13
rect 1782 -413 1803 -383
rect 291 -490 311 -450
rect 1728 -490 1748 -450
<< mvnsubdiff >>
rect 291 1251 311 1291
rect 1728 1251 1748 1291
rect 236 1194 257 1224
rect 0 485 20 525
rect 167 485 187 525
rect -54 425 -37 445
rect -54 145 -37 165
rect 236 140 257 157
rect 1782 1194 1803 1224
rect 1782 140 1803 157
<< mvpsubdiffcont >>
rect -54 -289 -37 -29
rect 236 -383 257 -30
rect 1782 -383 1803 -30
rect 311 -490 1728 -450
<< mvnsubdiffcont >>
rect 311 1251 1728 1291
rect 20 485 167 525
rect -54 165 -37 425
rect 236 157 257 1194
rect 1782 157 1803 1194
<< poly >>
rect 323 1224 373 1237
rect 402 1224 452 1237
rect 481 1224 531 1237
rect 560 1224 610 1237
rect 639 1224 689 1237
rect 718 1224 768 1237
rect 797 1224 847 1237
rect 876 1224 926 1237
rect 955 1224 1005 1237
rect 1034 1224 1084 1237
rect 1113 1224 1163 1237
rect 1192 1224 1242 1237
rect 1271 1224 1321 1237
rect 1350 1224 1400 1237
rect 1429 1224 1479 1237
rect 1508 1224 1558 1237
rect 1587 1224 1637 1237
rect 1666 1224 1716 1237
rect 29 445 79 458
rect 108 445 158 458
rect 29 116 79 145
rect 29 86 39 116
rect 69 86 79 116
rect 29 76 79 86
rect 108 116 158 145
rect 108 86 118 116
rect 148 86 158 116
rect 108 76 158 86
rect 323 60 373 140
rect 311 50 373 60
rect 311 20 321 50
rect 351 20 373 50
rect 311 10 373 20
rect 29 -9 79 4
rect 108 -9 158 4
rect 323 -13 373 10
rect 402 60 452 140
rect 481 60 531 140
rect 402 50 531 60
rect 402 20 424 50
rect 509 20 531 50
rect 402 10 531 20
rect 402 -13 452 10
rect 481 -13 531 10
rect 560 60 610 140
rect 639 60 689 140
rect 560 50 689 60
rect 560 20 582 50
rect 667 20 689 50
rect 560 10 689 20
rect 560 -13 610 10
rect 639 -13 689 10
rect 718 60 768 140
rect 797 60 847 140
rect 718 50 847 60
rect 718 20 740 50
rect 825 20 847 50
rect 718 10 847 20
rect 718 -13 768 10
rect 797 -13 847 10
rect 876 60 926 140
rect 955 60 1005 140
rect 876 50 1005 60
rect 876 20 898 50
rect 983 20 1005 50
rect 876 10 1005 20
rect 876 -13 926 10
rect 955 -13 1005 10
rect 1034 60 1084 140
rect 1113 60 1163 140
rect 1034 50 1163 60
rect 1034 20 1056 50
rect 1141 20 1163 50
rect 1034 10 1163 20
rect 1034 -13 1084 10
rect 1113 -13 1163 10
rect 1192 60 1242 140
rect 1271 60 1321 140
rect 1192 50 1321 60
rect 1192 20 1214 50
rect 1299 20 1321 50
rect 1192 10 1321 20
rect 1192 -13 1242 10
rect 1271 -13 1321 10
rect 1350 60 1400 140
rect 1429 60 1479 140
rect 1350 50 1479 60
rect 1350 20 1372 50
rect 1457 20 1479 50
rect 1350 10 1479 20
rect 1350 -13 1400 10
rect 1429 -13 1479 10
rect 1508 60 1558 140
rect 1587 60 1637 140
rect 1508 50 1637 60
rect 1508 20 1530 50
rect 1615 20 1637 50
rect 1508 10 1637 20
rect 1508 -13 1558 10
rect 1587 -13 1637 10
rect 1666 60 1716 140
rect 1666 50 1728 60
rect 1666 20 1688 50
rect 1718 20 1728 50
rect 1666 10 1728 20
rect 1666 -13 1716 10
rect 29 -338 79 -309
rect 29 -368 39 -338
rect 69 -368 79 -338
rect 29 -378 79 -368
rect 108 -338 158 -309
rect 108 -368 118 -338
rect 148 -368 158 -338
rect 108 -378 158 -368
rect 323 -426 373 -413
rect 402 -426 452 -413
rect 481 -426 531 -413
rect 560 -426 610 -413
rect 639 -426 689 -413
rect 718 -426 768 -413
rect 797 -426 847 -413
rect 876 -426 926 -413
rect 955 -426 1005 -413
rect 1034 -426 1084 -413
rect 1113 -426 1163 -413
rect 1192 -426 1242 -413
rect 1271 -426 1321 -413
rect 1350 -426 1400 -413
rect 1429 -426 1479 -413
rect 1508 -426 1558 -413
rect 1587 -426 1637 -413
rect 1666 -426 1716 -413
<< polycont >>
rect 39 86 69 116
rect 118 86 148 116
rect 321 20 351 50
rect 424 20 509 50
rect 582 20 667 50
rect 740 20 825 50
rect 898 20 983 50
rect 1056 20 1141 50
rect 1214 20 1299 50
rect 1372 20 1457 50
rect 1530 20 1615 50
rect 1688 20 1718 50
rect 39 -368 69 -338
rect 118 -368 148 -338
<< locali >>
rect 291 1251 311 1291
rect 1728 1251 1748 1291
rect 236 1194 257 1224
rect 0 485 20 525
rect 167 485 187 525
rect -54 425 -37 445
rect -54 145 -37 165
rect 6 439 23 447
rect 6 143 23 151
rect 85 439 102 447
rect 85 143 102 151
rect 164 439 181 447
rect 164 143 181 151
rect 236 140 257 157
rect 300 1218 317 1226
rect 300 138 317 146
rect 379 1218 396 1226
rect 379 138 396 146
rect 458 1218 475 1226
rect 458 138 475 146
rect 537 1218 554 1226
rect 537 138 554 146
rect 616 1218 633 1226
rect 616 138 633 146
rect 695 1218 712 1226
rect 695 138 712 146
rect 774 1218 791 1226
rect 774 138 791 146
rect 853 1218 870 1226
rect 853 138 870 146
rect 932 1218 949 1226
rect 932 138 949 146
rect 1011 1218 1028 1226
rect 1011 138 1028 146
rect 1090 1218 1107 1226
rect 1090 138 1107 146
rect 1169 1218 1186 1226
rect 1169 138 1186 146
rect 1248 1218 1265 1226
rect 1248 138 1265 146
rect 1327 1218 1344 1226
rect 1327 138 1344 146
rect 1406 1218 1423 1226
rect 1406 138 1423 146
rect 1485 1218 1502 1226
rect 1485 138 1502 146
rect 1564 1218 1581 1226
rect 1564 138 1581 146
rect 1643 1218 1660 1226
rect 1643 138 1660 146
rect 1722 1218 1739 1226
rect 1722 138 1739 146
rect 1782 1194 1803 1224
rect 1782 140 1803 157
rect 29 116 79 126
rect 29 86 39 116
rect 69 86 79 116
rect 29 60 79 86
rect 97 116 158 126
rect 97 86 107 116
rect 148 86 158 116
rect 97 76 158 86
rect 29 50 90 60
rect 29 20 50 50
rect 80 20 90 50
rect 29 10 90 20
rect 311 50 361 60
rect 311 20 321 50
rect 351 20 361 50
rect 311 10 361 20
rect 414 50 519 60
rect 414 20 424 50
rect 509 20 519 50
rect 414 10 519 20
rect 572 50 677 60
rect 572 20 582 50
rect 667 20 677 50
rect 572 10 677 20
rect 730 50 835 60
rect 730 20 740 50
rect 825 20 835 50
rect 730 10 835 20
rect 888 50 993 60
rect 888 20 898 50
rect 983 20 993 50
rect 888 10 993 20
rect 1046 50 1151 60
rect 1046 20 1056 50
rect 1141 20 1151 50
rect 1046 10 1151 20
rect 1204 50 1309 60
rect 1204 20 1214 50
rect 1299 20 1309 50
rect 1204 10 1309 20
rect 1362 50 1467 60
rect 1362 20 1372 50
rect 1457 20 1467 50
rect 1362 10 1467 20
rect 1520 50 1625 60
rect 1520 20 1530 50
rect 1615 20 1625 50
rect 1520 10 1625 20
rect 1678 50 1728 60
rect 1678 20 1688 50
rect 1718 20 1728 50
rect 1678 10 1728 20
rect -54 -29 -37 -9
rect -54 -309 -37 -289
rect 6 -15 23 -7
rect 6 -311 23 -303
rect 85 -15 102 -7
rect 85 -311 102 -303
rect 164 -15 181 -7
rect 164 -311 181 -303
rect 236 -30 257 -13
rect 29 -338 79 -328
rect 29 -368 39 -338
rect 69 -368 79 -338
rect 29 -489 79 -368
rect 108 -338 158 -328
rect 108 -368 118 -338
rect 148 -368 158 -338
rect 108 -489 158 -368
rect 236 -413 257 -383
rect 300 -19 317 -11
rect 300 -415 317 -407
rect 379 -19 396 -11
rect 379 -415 396 -407
rect 458 -19 475 -11
rect 458 -415 475 -407
rect 537 -19 554 -11
rect 537 -415 554 -407
rect 616 -19 633 -11
rect 616 -415 633 -407
rect 695 -19 712 -11
rect 695 -415 712 -407
rect 774 -19 791 -11
rect 774 -415 791 -407
rect 853 -19 870 -11
rect 853 -415 870 -407
rect 932 -19 949 -11
rect 932 -415 949 -407
rect 1011 -19 1028 -11
rect 1011 -415 1028 -407
rect 1090 -19 1107 -11
rect 1090 -415 1107 -407
rect 1169 -19 1186 -11
rect 1169 -415 1186 -407
rect 1248 -19 1265 -11
rect 1248 -415 1265 -407
rect 1327 -19 1344 -11
rect 1327 -415 1344 -407
rect 1406 -19 1423 -11
rect 1406 -415 1423 -407
rect 1485 -19 1502 -11
rect 1485 -415 1502 -407
rect 1564 -19 1581 -11
rect 1564 -415 1581 -407
rect 1643 -19 1660 -11
rect 1643 -415 1660 -407
rect 1722 -19 1739 -11
rect 1722 -415 1739 -407
rect 1782 -30 1803 -13
rect 1782 -413 1803 -383
rect 291 -490 311 -450
rect 1728 -490 1748 -450
<< viali >>
rect 311 1251 1728 1291
rect 20 485 167 525
rect -54 165 -37 425
rect 6 151 23 439
rect 85 151 102 439
rect 164 151 181 439
rect 236 157 257 1194
rect 300 146 317 1218
rect 379 146 396 1218
rect 458 146 475 1218
rect 537 146 554 1218
rect 616 146 633 1218
rect 695 146 712 1218
rect 774 146 791 1218
rect 853 146 870 1218
rect 932 146 949 1218
rect 1011 146 1028 1218
rect 1090 146 1107 1218
rect 1169 146 1186 1218
rect 1248 146 1265 1218
rect 1327 146 1344 1218
rect 1406 146 1423 1218
rect 1485 146 1502 1218
rect 1564 146 1581 1218
rect 1643 146 1660 1218
rect 1722 146 1739 1218
rect 1782 157 1803 1194
rect 107 86 118 116
rect 118 86 137 116
rect 50 20 80 50
rect 321 20 351 50
rect 424 20 509 50
rect 582 20 667 50
rect 740 20 825 50
rect 898 20 983 50
rect 1056 20 1141 50
rect 1214 20 1299 50
rect 1372 20 1457 50
rect 1530 20 1615 50
rect 1688 20 1718 50
rect -54 -289 -37 -29
rect 6 -303 23 -15
rect 85 -303 102 -15
rect 164 -303 181 -15
rect 236 -383 257 -30
rect 300 -407 317 -19
rect 379 -407 396 -19
rect 458 -407 475 -19
rect 537 -407 554 -19
rect 616 -407 633 -19
rect 695 -407 712 -19
rect 774 -407 791 -19
rect 853 -407 870 -19
rect 932 -407 949 -19
rect 1011 -407 1028 -19
rect 1090 -407 1107 -19
rect 1169 -407 1186 -19
rect 1248 -407 1265 -19
rect 1327 -407 1344 -19
rect 1406 -407 1423 -19
rect 1485 -407 1502 -19
rect 1564 -407 1581 -19
rect 1643 -407 1660 -19
rect 1722 -407 1739 -19
rect 1782 -383 1803 -30
rect 311 -490 1728 -450
<< metal1 >>
rect 226 1291 1813 1301
rect 226 1251 311 1291
rect 1728 1251 1813 1291
rect 226 1241 1813 1251
rect 226 1218 320 1241
rect 226 1194 300 1218
rect 226 535 236 1194
rect -64 525 236 535
rect -64 485 20 525
rect 167 485 236 525
rect -64 475 236 485
rect -64 425 -27 475
rect -64 165 -54 425
rect -37 165 -27 425
rect -64 145 -27 165
rect 3 439 26 445
rect 3 151 6 439
rect 23 151 26 439
rect 3 126 26 151
rect 82 439 105 475
rect 82 151 85 439
rect 102 151 105 439
rect 82 145 105 151
rect 161 439 184 445
rect 161 151 164 439
rect 181 151 184 439
rect 3 116 147 126
rect 3 86 107 116
rect 137 86 147 116
rect 3 76 147 86
rect -64 -29 -27 -9
rect -64 -289 -54 -29
rect -37 -289 -27 -29
rect -64 -349 -27 -289
rect 3 -15 26 76
rect 161 60 184 151
rect 226 157 236 475
rect 257 157 300 1194
rect 226 146 300 157
rect 317 146 320 1218
rect 226 140 320 146
rect 376 1218 399 1224
rect 376 146 379 1218
rect 396 146 399 1218
rect 376 125 399 146
rect 455 1218 478 1241
rect 455 146 458 1218
rect 475 146 478 1218
rect 455 140 478 146
rect 534 1218 557 1224
rect 534 146 537 1218
rect 554 146 557 1218
rect 534 125 557 146
rect 613 1218 636 1241
rect 613 146 616 1218
rect 633 146 636 1218
rect 613 140 636 146
rect 692 1218 715 1224
rect 692 146 695 1218
rect 712 146 715 1218
rect 692 125 715 146
rect 771 1218 794 1241
rect 771 146 774 1218
rect 791 146 794 1218
rect 771 140 794 146
rect 850 1218 873 1224
rect 850 146 853 1218
rect 870 146 873 1218
rect 850 125 873 146
rect 929 1218 952 1241
rect 929 146 932 1218
rect 949 146 952 1218
rect 929 140 952 146
rect 1008 1218 1031 1224
rect 1008 146 1011 1218
rect 1028 146 1031 1218
rect 1008 125 1031 146
rect 1087 1218 1110 1241
rect 1087 146 1090 1218
rect 1107 146 1110 1218
rect 1087 140 1110 146
rect 1166 1218 1189 1224
rect 1166 146 1169 1218
rect 1186 146 1189 1218
rect 1166 125 1189 146
rect 1245 1218 1268 1241
rect 1245 146 1248 1218
rect 1265 146 1268 1218
rect 1245 140 1268 146
rect 1324 1218 1347 1224
rect 1324 146 1327 1218
rect 1344 146 1347 1218
rect 1324 125 1347 146
rect 1403 1218 1426 1241
rect 1403 146 1406 1218
rect 1423 146 1426 1218
rect 1403 140 1426 146
rect 1482 1218 1505 1224
rect 1482 146 1485 1218
rect 1502 146 1505 1218
rect 1482 125 1505 146
rect 1561 1218 1584 1241
rect 1561 146 1564 1218
rect 1581 146 1584 1218
rect 1561 140 1584 146
rect 1640 1218 1663 1224
rect 1640 146 1643 1218
rect 1660 146 1663 1218
rect 1640 125 1663 146
rect 1719 1218 1813 1241
rect 1719 146 1722 1218
rect 1739 1194 1813 1218
rect 1739 157 1782 1194
rect 1803 157 1813 1194
rect 1739 146 1813 157
rect 1719 140 1813 146
rect 376 115 1728 125
rect 376 85 386 115
rect 1718 85 1728 115
rect 376 75 1728 85
rect 40 50 184 60
rect 40 20 50 50
rect 80 20 147 50
rect 177 20 184 50
rect 40 10 184 20
rect 311 50 361 60
rect 311 20 321 50
rect 351 20 361 50
rect 311 10 361 20
rect 3 -303 6 -15
rect 23 -303 26 -15
rect 3 -309 26 -303
rect 82 -15 105 -9
rect 82 -303 85 -15
rect 102 -303 105 -15
rect 82 -349 105 -303
rect 161 -15 184 10
rect 161 -303 164 -15
rect 181 -303 184 -15
rect 161 -309 184 -303
rect 226 -19 320 -13
rect 226 -30 300 -19
rect 226 -349 236 -30
rect -64 -383 236 -349
rect 257 -383 300 -30
rect -64 -407 300 -383
rect 317 -407 320 -19
rect -64 -409 320 -407
rect 226 -440 320 -409
rect 376 -19 399 75
rect 414 50 519 60
rect 414 20 424 50
rect 509 20 519 50
rect 414 10 519 20
rect 376 -407 379 -19
rect 396 -407 399 -19
rect 376 -413 399 -407
rect 455 -19 478 -13
rect 455 -407 458 -19
rect 475 -407 478 -19
rect 455 -440 478 -407
rect 534 -19 557 75
rect 572 50 677 60
rect 572 20 582 50
rect 667 20 677 50
rect 572 10 677 20
rect 534 -407 537 -19
rect 554 -407 557 -19
rect 534 -413 557 -407
rect 613 -19 636 -13
rect 613 -407 616 -19
rect 633 -407 636 -19
rect 613 -440 636 -407
rect 692 -19 715 75
rect 730 50 835 60
rect 730 20 740 50
rect 825 20 835 50
rect 730 10 835 20
rect 692 -407 695 -19
rect 712 -407 715 -19
rect 692 -413 715 -407
rect 771 -19 794 -13
rect 771 -407 774 -19
rect 791 -407 794 -19
rect 771 -440 794 -407
rect 850 -19 873 75
rect 888 50 993 60
rect 888 20 898 50
rect 983 20 993 50
rect 888 10 993 20
rect 850 -407 853 -19
rect 870 -407 873 -19
rect 850 -413 873 -407
rect 929 -19 952 -13
rect 929 -407 932 -19
rect 949 -407 952 -19
rect 929 -440 952 -407
rect 1008 -19 1031 75
rect 1046 50 1151 60
rect 1046 20 1056 50
rect 1141 20 1151 50
rect 1046 10 1151 20
rect 1008 -407 1011 -19
rect 1028 -407 1031 -19
rect 1008 -413 1031 -407
rect 1087 -19 1110 -13
rect 1087 -407 1090 -19
rect 1107 -407 1110 -19
rect 1087 -440 1110 -407
rect 1166 -19 1189 75
rect 1204 50 1309 60
rect 1204 20 1214 50
rect 1299 20 1309 50
rect 1204 10 1309 20
rect 1166 -407 1169 -19
rect 1186 -407 1189 -19
rect 1166 -413 1189 -407
rect 1245 -19 1268 -13
rect 1245 -407 1248 -19
rect 1265 -407 1268 -19
rect 1245 -440 1268 -407
rect 1324 -19 1347 75
rect 1362 50 1467 60
rect 1362 20 1372 50
rect 1457 20 1467 50
rect 1362 10 1467 20
rect 1324 -407 1327 -19
rect 1344 -407 1347 -19
rect 1324 -413 1347 -407
rect 1403 -19 1426 -13
rect 1403 -407 1406 -19
rect 1423 -407 1426 -19
rect 1403 -440 1426 -407
rect 1482 -19 1505 75
rect 1520 50 1625 60
rect 1520 20 1530 50
rect 1615 20 1625 50
rect 1520 10 1625 20
rect 1482 -407 1485 -19
rect 1502 -407 1505 -19
rect 1482 -413 1505 -407
rect 1561 -19 1584 -13
rect 1561 -407 1564 -19
rect 1581 -407 1584 -19
rect 1561 -440 1584 -407
rect 1640 -19 1663 75
rect 1678 50 1728 60
rect 1678 20 1688 50
rect 1718 20 1728 50
rect 1678 10 1728 20
rect 1640 -407 1643 -19
rect 1660 -407 1663 -19
rect 1640 -413 1663 -407
rect 1719 -19 1813 -13
rect 1719 -407 1722 -19
rect 1739 -30 1813 -19
rect 1739 -383 1782 -30
rect 1803 -383 1813 -30
rect 1739 -407 1813 -383
rect 1719 -440 1813 -407
rect 226 -450 1813 -440
rect 226 -490 311 -450
rect 1728 -490 1813 -450
rect 226 -500 1813 -490
<< via1 >>
rect 386 85 1718 115
rect 147 20 177 50
rect 321 20 351 50
rect 424 20 509 50
rect 582 20 667 50
rect 740 20 825 50
rect 898 20 983 50
rect 1056 20 1141 50
rect 1214 20 1299 50
rect 1372 20 1457 50
rect 1530 20 1615 50
rect 1688 20 1718 50
<< metal2 >>
rect 376 115 1836 125
rect 376 85 386 115
rect 1718 85 1836 115
rect 376 75 1836 85
rect 137 50 1728 60
rect 137 20 147 50
rect 177 20 321 50
rect 351 20 424 50
rect 509 20 582 50
rect 667 20 740 50
rect 825 20 898 50
rect 983 20 1056 50
rect 1141 20 1214 50
rect 1299 20 1372 50
rect 1457 20 1530 50
rect 1615 20 1688 50
rect 1718 20 1728 50
rect 137 10 1728 20
<< labels >>
rlabel locali 29 -489 79 -439 5 Q
rlabel locali 108 -489 158 -439 5 QN
rlabel metal2 1786 75 1836 125 3 out
rlabel metal1 231 1251 281 1301 1 VH
rlabel metal1 231 -500 281 -450 5 VL
<< end >>
