* NGSPICE file created from converter_3.ext - technology: sky130A

.subckt level_shifter level_shifter_0/GND level_shifter_0/OUT
X0 a_1660_2346# level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X1 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X2 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X3 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X4 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X5 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X6 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X7 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X8 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X9 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X10 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X11 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X12 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X13 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.6 as=2.9 ps=20.3 w=20 l=0.5
X14 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X15 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X16 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X17 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X18 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X19 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X20 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/VDD level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X21 level_shifter_0/cruzados_0/OUT level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X22 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X23 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X24 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X25 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/VDD level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X26 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X27 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X28 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X29 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X30 level_shifter_0/VDD level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X31 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X32 level_shifter_0/cruzados_0/OUT a_1660_2346# level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X33 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X34 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=5.8 ps=40.6 w=20 l=0.5
X35 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X36 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=0.5
X37 level_shifter_0/cruzados_0/OUT level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X38 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X39 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X40 level_shifter_0/GND level_shifter_0/IN a_1660_2346# level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X41 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X42 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=5.8 ps=40.6 w=20 l=0.5
X43 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X44 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X45 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X46 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X47 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X48 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/VDD level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X49 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X50 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X51 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=0.5
X52 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X53 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=0.5
X54 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X55 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X56 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X57 level_shifter_0/GND level_shifter_0/inv_1_8_0/OUT level_shifter_0/cruzados_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X58 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X59 a_1660_2346# level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X60 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=5.8 pd=40.6 as=2.9 ps=20.3 w=20 l=0.5
X61 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X62 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X63 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X64 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=0.5
X65 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X66 level_shifter_0/VDD level_shifter_0/IN level_shifter_0/inv_1_8_0/OUT level_shifter_0/VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X67 level_shifter_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X68 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X69 level_shifter_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X70 level_shifter_0/GND level_shifter_0/IN level_shifter_0/inv_400_0/IN level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X71 level_shifter_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X72 level_shifter_0/inv_1_8_0/OUT level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X73 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
X74 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/VH level_shifter_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X75 level_shifter_0/inv_400_0/IN level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X76 a_1660_2346# level_shifter_0/IN level_shifter_0/GND level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X77 level_shifter_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/OUT level_shifter_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=0.5
.ends

.subckt nmos_drain_in m5_0_0# m4_648_1020# a_n6_62# dw_0_0# m3_0_0# w_0_0# a_100_62#
+ m5_788_894# m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.78 ps=18.8 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=2.78 pd=18.8 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_source_in m5_0_0# m4_648_1020# a_n6_62# dw_0_0# m3_0_0# w_0_0# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# w_0_0# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.86 ps=16.6 w=4.38 l=0.5
X1 w_0_0# a_0_0# a_n6_62# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=6.86 pd=16.6 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_source_frame_lt m4_n1950_0# m4_648_1020# m5_n1950_0# a_n950_0# m5_788_894#
+ m3_n1950_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_n950_0# a_n950_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=12.5 ps=32.6 w=4.38 l=0.5
.ends

.subckt nmos_drain_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020# a_1550_0#
X0 a_162_1100# a_0_0# a_100_62# a_1550_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=2.03 ps=14.1 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# a_1550_0# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.1 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_source_frame_rb m5_0_0# m4_648_1020# a_n6_62# m3_0_0# a_100_62# m5_788_894#
+ m4_0_0# a_0_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_100_62# a_100_62# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=6.23 ps=16.3 w=4.38 l=0.5
X1 a_100_62# a_0_0# a_n6_62# a_100_62# sky130_fd_pr__nfet_g5v0d10v5 ad=6.23 pd=16.3 as=0.131 ps=8.82 w=4.38 l=0.5
.ends

.subckt nmos_drain_frame_lt m4_648_1020# m3_n950_0# a_n950_0# m4_n950_0# m5_n950_0#
+ m5_788_894# a_0_0# a_162_0# a_162_1100# m3_648_1020#
X0 a_162_1100# a_0_0# a_162_0# a_n950_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=4.05 ps=28.2 w=4.38 l=0.5
.ends

.subckt nmos_waffle_36x36 a_n938_0# a_37562_0# a_n1100_n1200#
Xnmos_drain_in_574 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_541 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_552 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_530 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_563 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_305 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_338 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_316 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_349 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_327 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_135 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_168 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_371 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_113 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_146 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_382 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_179 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_124 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_102 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_360 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_393 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_157 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_28 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_17 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_39 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_190 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_8 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_509 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_520 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_531 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_339 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_542 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_575 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_317 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_553 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_328 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_306 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_564 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_372 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_383 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_350 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_103 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_394 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_361 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_169 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_147 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_114 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_125 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_158 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_136 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_29 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_18 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_180 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_191 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_9 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_543 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_576 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_521 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_318 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_554 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_329 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_532 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_565 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_307 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_510 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_373 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_351 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_384 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_362 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_340 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_395 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_115 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_148 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_159 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_126 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_137 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_104 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_19 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_181 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_192 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_170 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_490 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_577 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_522 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_319 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_555 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_500 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_566 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_533 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_511 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_544 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_308 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_352 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_149 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_116 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_385 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_127 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_330 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_396 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_363 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_341 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_374 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_105 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_138 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_182 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_160 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_193 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_171 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_491 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_480 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_556 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_523 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_501 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_534 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_567 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_545 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_309 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_512 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_320 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_117 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_386 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_353 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_128 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_331 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_364 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_397 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_375 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_139 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_342 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_106 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_30 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_150 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_183 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_161 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_172 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_194 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_492 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_470 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_481 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_524 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_557 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_535 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_502 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_568 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_546 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_513 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_0 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_118 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_354 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_321 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_387 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_129 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_365 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_332 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_398 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_107 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_376 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_310 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_343 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_20 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_184 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_151 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_31 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_195 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_162 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_140 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_173 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_471 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_482 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_460 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_493 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_290 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_525 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_503 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_536 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_547 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_514 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_558 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_569 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_30 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_322 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_388 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_355 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_300 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_333 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_399 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_366 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_311 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_108 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_119 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_1 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_344 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_377 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_32 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_lt_10 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_152 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_185 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_130 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_163 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_21 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_196 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_141 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_174 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_472 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_450 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_483 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_494 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_461 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_280 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_291 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_526 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_559 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_504 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_537 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_515 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_548 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_20 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_31 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_356 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_389 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_334 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_301 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_367 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_312 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_345 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_323 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_2 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_378 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_109 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_frame_lt_22 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_186 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_33 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_164 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_131 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_197 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_142 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_175 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_11 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_120 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_153 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_473 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_440 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_484 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_451 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_495 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_462 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_270 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_281 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_292 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_538 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_505 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_516 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_549 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_527 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_32 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_10 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_21 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_302 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_313 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_3 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_368 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_335 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_346 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_379 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_357 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_324 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_12 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_132 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_198 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_165 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_23 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_110 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_176 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_143 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_187 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_154 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_121 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_430 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_441 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_474 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_452 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_485 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_463 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_496 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_271 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_282 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_260 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_293 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_506 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_539 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_517 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_528 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_22 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_33 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_11 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_4 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_336 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_303 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_369 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_314 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_347 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_358 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_325 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_24 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_100 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_133 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_166 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_111 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_144 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_177 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_13 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_188 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_122 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_155 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_199 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_475 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_453 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_420 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_486 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_431 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_464 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_442 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_497 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_283 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_250 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_261 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_294 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_272 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_507 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_518 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_529 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_12 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_23 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_5 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_304 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_337 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_315 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_348 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_326 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_359 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_14 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_101 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_134 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_167 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_25 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_145 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_112 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_178 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_156 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_189 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_123 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_421 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_487 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_454 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_465 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_432 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_498 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_476 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_443 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_410 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_251 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_284 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_295 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_262 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_273 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_240 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_508 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_519 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_24 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_13 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_305 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_338 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_349 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_316 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_6 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_0 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_327 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_26 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_135 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_168 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_113 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_179 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_146 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_15 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_124 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_102 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_157 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_455 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_422 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_488 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_400 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_433 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_499 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_466 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_477 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_411 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_444 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_285 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_252 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_230 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_263 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_296 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_241 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_274 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_509 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_14 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_25 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_339 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_1 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_317 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_328 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_7 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_306 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_16 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_169 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_114 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_27 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_147 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_158 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_125 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_136 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_103 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_423 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_456 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_489 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_401 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_434 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_467 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_445 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_478 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_412 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_220 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_253 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_286 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_264 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_231 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_297 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_275 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_242 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_90 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_26 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_15 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_318 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_329 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_2 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_rb_8 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_307 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_28 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_148 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_115 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_17 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_126 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_159 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_137 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_104 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_424 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_402 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_435 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_413 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_446 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_457 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_468 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_479 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_254 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_490 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_287 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_232 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_298 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_265 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_243 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_210 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_221 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_276 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_0 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_80 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_91 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_16 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_27 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_rb_9 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_lt_3 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_319 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_308 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_18 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_116 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_29 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_149 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_127 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_138 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_105 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_458 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_403 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_436 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_469 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_447 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_414 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_425 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_288 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_491 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_233 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_200 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_266 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_299 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_211 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_277 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_244 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_222 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_255 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_480 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_1 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_81 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_92 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_70 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_28 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_17 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_4 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_309 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_117 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_19 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_in_128 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_106 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_139 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_404 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_437 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_415 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_448 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_426 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_459 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_492 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_201 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_470 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_212 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_481 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_234 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_267 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_245 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_278 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_256 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_289 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_2 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_223 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_82 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_93 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_60 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_71 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_18 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_rb_29 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_5 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_118 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_129 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_107 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_405 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_438 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_416 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_449 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_427 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_471 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_482 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_493 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_460 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_235 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_202 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_268 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_246 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_213 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_279 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_257 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_3 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_224 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_290 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_50 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_83 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_61 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_94 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_72 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_19 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_6 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_in_108 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_119 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_406 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_439 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_417 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_428 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_203 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_269 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_236 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_472 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_214 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_450 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_247 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_483 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_494 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_461 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_225 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_258 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_4 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_280 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_291 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_84 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_62 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_95 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_40 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_73 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_51 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_7 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_0 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_in_109 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_407 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_418 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_429 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_237 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_440 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_473 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_215 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_451 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_248 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_484 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_226 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_204 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_462 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_495 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_259 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_5 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_270 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_281 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_292 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_30 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_96 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_63 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_74 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_41 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_52 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_85 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_rb_1 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_drain_frame_lt_8 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_in_419 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_408 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_441 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_474 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_249 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_216 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_485 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_452 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_227 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_430 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_238 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_205 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_496 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_463 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_6 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_271 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_282 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_260 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_293 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_31 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_64 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_97 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_42 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_75 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_86 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_20 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_53 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_9 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_2 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_409 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_475 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_420 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_217 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_453 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_486 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_228 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_464 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_431 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_442 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_206 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_497 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_7 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_239 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_250 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_283 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_294 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_261 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_272 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_32 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_98 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_65 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_570 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_43 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_10 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_76 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_54 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_87 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_21 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_lt_30 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_3 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_90 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_454 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_421 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_487 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_432 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_498 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_465 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_443 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_476 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_410 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_218 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_229 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_8 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_207 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_284 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_251 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_262 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_295 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_273 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_240 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_560 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_33 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_11 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_571 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_44 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_22 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_55 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_66 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_99 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_77 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_88 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_390 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_31 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_20 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_4 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_80 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_91 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_422 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_400 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_411 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_219 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_455 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_488 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_433 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_466 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_499 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_477 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_444 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_208 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_9 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_252 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_285 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_263 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_230 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_296 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_274 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_241 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_30 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_67 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_12 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_572 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_45 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_78 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_550 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_56 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_23 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_34 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_561 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_89 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_380 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_391 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_21 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_32 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_10 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_5 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_81 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_92 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_70 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_456 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_423 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_489 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_401 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_467 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_434 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_209 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_478 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_412 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_445 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_220 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_286 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_253 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_231 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_297 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_264 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_242 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_275 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_31 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_20 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_573 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_540 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_46 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_13 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_79 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_551 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_24 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_57 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_68 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_35 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_562 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_370 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_381 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_392 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_33 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_11 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_22 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_6 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_0 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_82 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_60 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_93 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_71 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_424 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_457 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_402 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_435 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_468 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_413 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_446 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_479 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_254 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_287 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_232 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_21 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_265 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_298 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_210 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_243 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_32 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_221 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_10 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_276 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_541 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_14 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_574 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_47 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_552 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_25 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_58 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_69 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_36 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_563 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_530 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_371 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_382 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_393 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_360 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_23 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_12 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_1 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_frame_rb_7 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_190 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_50 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_83 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_94 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_61 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_72 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_458 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_403 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_436 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_469 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_414 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_447 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_425 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_288 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_200 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_266 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_233 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_299 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_244 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_211 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_277 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_255 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_222 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_33 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_575 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_542 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_48 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_15 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_520 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_553 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_59 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_26 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_11 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_564 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_531 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_22 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_37 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_372 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_350 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_383 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_361 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_394 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_13 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_2 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_frame_lt_24 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_8 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_in_180 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_191 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_84 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_62 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_95 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_73 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_40 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_51 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_404 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_437 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_448 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_415 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_459 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_426 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_234 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_201 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_267 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_212 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_278 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_245 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_289 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_256 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_223 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_543 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_16 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_576 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_49 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_23 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_521 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_554 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_27 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_532 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_565 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_510 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_12 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_38 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_373 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_351 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_384 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_362 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_340 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_395 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_25 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_14 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_rb_9 a_n938_0# a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0#
+ a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_rb
Xnmos_source_frame_lt_3 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_181 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_192 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_170 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_30 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_63 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_96 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_41 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_74 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_85 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_52 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_405 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_438 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_416 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_427 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_449 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_202 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_235 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_268 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_213 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_246 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_279 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_224 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_257 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_555 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_522 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_13 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_533 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_500 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_544 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_24 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_511 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_577 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_28 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_566 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_39 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_17 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_385 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_352 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_363 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_330 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_396 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_374 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_341 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_15 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_26 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_4 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_182 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_193 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_160 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_171 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_31 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_97 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_64 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_42 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_75 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_86 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_53 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_20 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_406 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_439 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_417 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_428 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_0 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_203 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_236 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_269 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_247 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_214 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_258 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_225 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_25 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_frame_rb_14 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_523 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_556 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_29 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_501 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_567 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_534 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_18 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_545 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_512 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_353 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_320 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_386 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_331 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_397 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_364 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_375 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_342 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_27 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_16 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_5 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_183 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_150 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_161 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_194 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_172 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_65 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_32 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_98 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_10 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_76 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_43 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_87 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_21 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_54 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_407 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_418 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_429 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_1 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_204 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_237 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_215 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_248 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_15 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_226 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_26 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_drain_in_259 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_557 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_524 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_502 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_535 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_568 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_19 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_513 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_546 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_321 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_310 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_387 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_354 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_332 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_365 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_398 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_343 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_376 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_17 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_6 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_drain_frame_lt_28 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_in_151 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_184 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_162 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_195 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_173 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_140 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_33 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_99 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_66 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_11 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_44 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_77 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_22 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_55 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_88 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_419 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_408 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_2 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_216 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_249 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_227 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_205 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_238 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_525 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_558 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_27 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_536 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_503 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_569 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_16 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_547 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_514 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_322 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_355 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_388 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_300 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_366 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_333 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_399 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_311 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_377 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_344 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_29 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_drain_frame_lt_18 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_7 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_152 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_185 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_130 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_196 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_163 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_141 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_174 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_12 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_67 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_45 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_78 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_23 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_56 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_34 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_89 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_409 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_3 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_217 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_228 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_239 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_206 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_526 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_559 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_504 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_537 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_17 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_515 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_548 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_28 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_356 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_389 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_301 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_334 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_367 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_570 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_345 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_312 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_323 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_378 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_lt_19 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_37562_0#
+ a_n1100_n1200# a_n938_0# a_37562_0# a_37562_0# nmos_drain_frame_lt
Xnmos_source_frame_lt_8 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_186 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_131 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_164 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_197 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_175 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_142 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_120 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_153 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_13 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_79 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_46 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_57 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_24 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_35 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_68 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_4 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_218 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_229 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_207 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_29 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_505 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_538 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_549 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_516 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_frame_rb_18 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_527 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_560 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_335 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_302 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_368 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_571 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_313 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_379 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_346 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_324 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_357 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_390 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_frame_lt_9 a_n938_0# a_n938_0# a_n938_0# a_37562_0# a_n938_0# a_n938_0#
+ a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_frame_lt
Xnmos_source_in_132 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_165 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_198 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_110 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_143 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_176 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_154 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_187 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_121 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_47 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_14 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_25 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_58 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_69 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_36 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_5 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_219 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_208 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_frame_rb_19 a_37562_0# a_37562_0# a_37562_0# a_37562_0# a_n938_0# a_37562_0#
+ a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# a_37562_0# nmos_drain_frame_rb
Xnmos_source_in_506 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_539 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_517 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_528 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_303 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_336 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_369 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_572 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_314 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_550 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_347 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_561 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_358 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_325 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_133 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_100 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_199 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_166 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_144 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_111 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_380 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_177 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_391 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_188 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_155 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_122 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_15 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_48 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_26 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_59 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_37 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_6 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_209 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_507 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_518 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_529 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_337 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_304 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_540 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_573 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_315 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_551 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_562 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_326 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_348 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_359 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_101 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_167 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_134 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_370 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_112 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_178 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_145 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_drain_in_381 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_drain_in_392 a_37562_0# a_37562_0# a_37562_0# dw_n6950_n7050# a_37562_0# a_37562_0#
+ a_n938_0# a_37562_0# a_37562_0# a_n1100_n1200# a_37562_0# a_37562_0# nmos_drain_in
Xnmos_source_in_189 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_123 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_156 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_16 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_49 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_27 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_38 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_7 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_508 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
Xnmos_source_in_519 a_n938_0# a_n938_0# a_n938_0# dw_n6950_n7050# a_n938_0# a_37562_0#
+ a_n938_0# a_n938_0# a_n1100_n1200# a_n938_0# a_n938_0# nmos_source_in
X0 a_37562_0# a_n1100_n1200# a_n938_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=1.33 ps=9.38 w=4.38 l=0.5
X1 a_37562_0# a_n1100_n1200# a_n938_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=11.2 pd=32 as=0.131 ps=8.82 w=4.38 l=0.5
X2 a_n938_0# a_n1100_n1200# a_37562_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=9.38 as=0.131 ps=8.82 w=4.38 l=0.5
X3 a_n938_0# a_n1100_n1200# a_37562_0# a_37562_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0.131 pd=8.82 as=11.2 ps=32 w=4.38 l=0.5
.ends

.subckt power_stage_3 VP out s2 VN
Xnmos_waffle_36x36_0 out VN s1 nmos_waffle_36x36
Xnmos_waffle_36x36_1 VP out s2 nmos_waffle_36x36
.ends

.subckt mimcap_30x30 c2_30_30# c1_30_30# m3_0_0#
X0 c1_30_30# m3_0_0# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X1 c2_30_30# c1_30_30# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt mimcap_210x420 mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0# mimcap_30x30_9/c2_30_30#
Xmimcap_30x30_90 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_80 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_91 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_70 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_81 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_92 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_60 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_71 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_82 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_93 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_50 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_61 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_72 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_83 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_94 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_40 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_51 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_62 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_73 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_84 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_95 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_96 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_30 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_41 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_52 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_63 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_74 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_85 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_97 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_20 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_31 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_42 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_53 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_64 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_75 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_86 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_21 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_10 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_32 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_43 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_54 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_65 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_76 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_87 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_22 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_11 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_0 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_33 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_44 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_55 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_66 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_77 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_88 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_23 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_12 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_34 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_45 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_56 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_67 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_78 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_89 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_1 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_2 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_24 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_13 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_35 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_46 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_57 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_68 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_79 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_14 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_25 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_36 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_47 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_58 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_69 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_3 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_15 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_4 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_26 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_37 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_48 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_59 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_16 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_27 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_38 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_49 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_5 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_17 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_28 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_39 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_6 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_18 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_29 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_7 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_19 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_8 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
Xmimcap_30x30_9 mimcap_30x30_9/c2_30_30# mimcap_30x30_9/c1_30_30# mimcap_30x30_9/m3_0_0#
+ mimcap_30x30
.ends

.subckt boot_ls_stage w_n1158_n782# RESET SET VDD GND
X0 VDD RESET RESET VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X1 w_n1158_n782# Iref GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X2 VDD RESET w_n1370_986# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 w_n1158_n782# VFE RESET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 GND Iref w_n1158_n782# GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=2
X5 w_n1158_n782# VRE SET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 RESET VFE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 RESET VFE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 SET SET VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X9 SET VRE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 SET SET w_n1370_986# w_n1370_986# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 w_888_986# RESET RESET w_888_986# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 w_n1158_n782# VRE SET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 w_n1158_n782# VFE RESET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 w_888_986# SET VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X15 GND Iref Iref GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=2
X16 VDD SET RESET VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=1
X17 SET VRE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X18 SET RESET VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=1
X19 w_n1158_n782# VRE SET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X20 w_n1158_n782# VFE RESET w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X21 SET VRE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X22 RESET VFE w_n1158_n782# w_n1158_n782# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt buffer QN Q VDD VSS
X0 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X1 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 VSS Q a_n195_154# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X4 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X7 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_n137_16# a_n195_154# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.475 ps=3.37 w=3 l=0.5
X10 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X11 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X12 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X13 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X14 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X15 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X16 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X17 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X18 VDD a_n137_16# a_n195_154# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.475 pd=3.37 as=0.29 ps=2.58 w=1 l=0.5
X19 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X20 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X21 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X22 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=3.14 ps=22.3 w=10.8 l=0.5
X23 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X24 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X25 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X26 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=3.14 pd=22.3 as=1.57 ps=11.1 w=10.8 l=0.5
X27 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X28 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X29 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X30 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X31 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X32 a_n137_16# QN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X33 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X34 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X35 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X36 out a_n137_16# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X37 out a_n137_16# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X38 VDD a_n137_16# out VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.57 pd=11.1 as=1.57 ps=11.1 w=10.8 l=0.5
X39 VSS a_n137_16# out VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt nand_5v B A AND VDD GND
X0 a_n29_n1168# B GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=3
X1 AND B VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=3
X2 AND A a_n29_n1168# GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=3
X3 VDD A AND VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=3
.ends

.subckt driver_bootstrap w_n3969_322# VBOOT VSUBS buffer_0/VSS
Xboot_ls_stage_0 w_n3969_322# nand_5v_1/A nand_5v_0/A VBOOT VSUBS boot_ls_stage
Xbuffer_0 nand_5v_1/B buffer_0/Q VBOOT buffer_0/VSS buffer
Xnand_5v_0 buffer_0/Q nand_5v_0/A nand_5v_1/B VBOOT buffer_0/VSS nand_5v
Xnand_5v_1 nand_5v_1/B nand_5v_1/A buffer_0/Q VBOOT buffer_0/VSS nand_5v
.ends

.subckt converter_3
Xlevel_shifter_0 VSUBS power_stage_3_0/s2 level_shifter
Xpower_stage_3_0 VSS Vout power_stage_3_0/s2 VDD power_stage_3
Xmimcap_210x420_0 driver_bootstrap_0/VBOOT Vout Vout mimcap_210x420
Xdriver_bootstrap_0 w_108020_n12608# driver_bootstrap_0/VBOOT VSUBS driver_bootstrap_0/buffer_0/VSS
+ driver_bootstrap
.ends

