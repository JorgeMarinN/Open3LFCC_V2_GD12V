magic
tech sky130A
magscale 1 2
timestamp 1699908495
<< metal2 >>
rect 10382 6360 10702 6400
rect 10382 5440 10422 6360
rect 10662 5440 10702 6360
rect 10382 -800 10702 5440
<< via2 >>
rect 10422 5440 10662 6360
<< metal3 >>
rect 10382 6360 10702 6400
rect 10382 5440 10422 6360
rect 10662 5440 10702 6360
rect 10382 -800 10702 5440
rect 18000 1560 104000 1600
rect 18000 440 18040 1560
rect 103960 440 104000 1560
rect 18000 0 104000 440
rect 106000 -2040 108000 -2000
rect 106000 -43960 106040 -2040
rect 107960 -43960 108000 -2040
rect 106000 -44000 108000 -43960
<< via3 >>
rect 10422 5440 10662 6360
rect 18040 440 103960 1560
rect 106040 -43960 107960 -2040
<< metal4 >>
rect 10382 6360 10702 6400
rect 10382 5440 10422 6360
rect 10662 5440 10702 6360
rect 10382 -800 10702 5440
rect 18000 1560 104000 2000
rect 18000 440 18040 1560
rect 103960 440 104000 1560
rect 18000 400 104000 440
rect 105320 -2040 108000 -2000
rect 105320 -43960 106040 -2040
rect 107960 -43960 108000 -2040
rect 105320 -44000 108000 -43960
<< via4 >>
rect 10422 5440 10662 6360
rect 18040 440 103960 1560
<< metal5 >>
rect 2000 56000 6000 60000
rect 116000 56000 120000 60000
rect 60000 46000 64000 50000
rect 10382 6360 10702 6400
rect 10382 5440 10422 6360
rect 10662 5440 10702 6360
rect 10382 -800 10702 5440
rect 18000 1560 104000 1600
rect 18000 440 18040 1560
rect 103960 440 104000 1560
rect 18000 0 104000 440
use driver_bootstrap  driver_bootstrap_0
timestamp 1699906343
transform 1 0 114255 0 1 -4348
box -4255 -1652 7801 2666
use level_shifter  level_shifter_0
timestamp 1699906343
transform 0 -1 14936 1 0 -6600
box 0 0 6050 8936
use mimcap_210x420  mimcap_210x420_0
timestamp 1699906343
transform 1 0 16000 0 1 -44660
box 0 0 89320 44660
use power_stage_3  power_stage_3_0
timestamp 1699906343
transform 0 1 0 1 0 0
box 0 0 61200 123200
<< labels >>
rlabel metal5 2000 56000 6000 60000 1 VSS
rlabel metal5 116000 56000 120000 60000 1 VDD
rlabel metal5 60000 46000 64000 50000 1 Vout
<< end >>
