magic
tech sky130A
magscale 1 2
timestamp 1698878589
<< dnwell >>
rect -1074 -1554 1074 106
<< nwell >>
rect -887 186 887 1368
rect -1154 -100 1154 186
rect -1154 -1348 -868 -100
rect 868 -1348 1154 -100
rect -1154 -1634 1154 -1348
<< pwell >>
rect -868 -1348 868 -100
<< mvnmos >>
rect -629 -1168 -29 -168
rect 29 -1168 629 -168
<< mvpmos >>
rect -629 168 -29 1168
rect 29 168 629 1168
<< mvndiff >>
rect -687 -180 -629 -168
rect -687 -1156 -675 -180
rect -641 -1156 -629 -180
rect -687 -1168 -629 -1156
rect -29 -180 29 -168
rect -29 -1156 -17 -180
rect 17 -1156 29 -180
rect -29 -1168 29 -1156
rect 629 -180 687 -168
rect 629 -1156 641 -180
rect 675 -1156 687 -180
rect 629 -1168 687 -1156
<< mvpdiff >>
rect -687 1156 -629 1168
rect -687 180 -675 1156
rect -641 180 -629 1156
rect -687 168 -629 180
rect -29 1156 29 1168
rect -29 180 -17 1156
rect 17 180 29 1156
rect -29 168 29 180
rect 629 1156 687 1168
rect 629 180 641 1156
rect 675 180 687 1156
rect 629 168 687 180
<< mvndiffc >>
rect -675 -1156 -641 -180
rect -17 -1156 17 -180
rect 641 -1156 675 -180
<< mvpdiffc >>
rect -675 180 -641 1156
rect -17 180 17 1156
rect 641 180 675 1156
<< mvpsubdiff >>
rect -841 -198 -761 -168
rect -841 -1138 -821 -198
rect -781 -1138 -761 -198
rect -841 -1168 -761 -1138
rect 761 -198 841 -168
rect 761 -1138 781 -198
rect 821 -1138 841 -198
rect 761 -1168 841 -1138
rect -687 -1262 687 -1242
rect -687 -1302 -657 -1262
rect 657 -1302 687 -1262
rect -687 -1322 687 -1302
<< mvnsubdiff >>
rect -687 1282 687 1302
rect -687 1242 -657 1282
rect 657 1242 687 1282
rect -687 1222 687 1242
rect -821 1138 -741 1168
rect -821 198 -801 1138
rect -761 198 -741 1138
rect -821 168 -741 198
rect 741 1138 821 1168
rect 741 198 761 1138
rect 801 198 821 1138
rect 741 168 821 198
rect -1074 -200 -994 -170
rect -1074 -1318 -1054 -200
rect -1014 -1318 -994 -200
rect 994 -200 1074 -170
rect -1074 -1348 -994 -1318
rect 994 -1318 1014 -200
rect 1054 -1318 1074 -200
rect 994 -1348 1074 -1318
rect -868 -1494 868 -1474
rect -868 -1534 -838 -1494
rect 838 -1534 868 -1494
rect -868 -1554 868 -1534
<< mvpsubdiffcont >>
rect -821 -1138 -781 -198
rect 781 -1138 821 -198
rect -657 -1302 657 -1262
<< mvnsubdiffcont >>
rect -657 1242 657 1282
rect -801 198 -761 1138
rect 761 198 801 1138
rect -1054 -1318 -1014 -200
rect 1014 -1318 1054 -200
rect -838 -1534 838 -1494
<< poly >>
rect -629 1168 -29 1194
rect 29 1168 629 1194
rect -629 142 -29 168
rect 29 142 629 168
rect -607 94 -51 142
rect -607 34 -587 94
rect -71 34 -51 94
rect -607 -142 -51 34
rect 51 -34 607 142
rect 51 -94 71 -34
rect 587 -94 607 -34
rect 51 -142 607 -94
rect -629 -168 -29 -142
rect 29 -168 629 -142
rect -629 -1194 -29 -1168
rect 29 -1194 629 -1168
<< polycont >>
rect -587 34 -71 94
rect 71 -94 587 -34
<< locali >>
rect -687 1282 687 1302
rect -687 1242 -657 1282
rect 657 1242 687 1282
rect -687 1222 687 1242
rect -821 1138 -741 1168
rect -821 300 -801 1138
rect -1074 200 -801 300
rect -1074 -200 -994 200
rect -821 198 -801 200
rect -761 198 -741 1138
rect -821 168 -741 198
rect -675 1156 -641 1172
rect -675 164 -641 180
rect -17 1156 17 1172
rect -17 164 17 180
rect 641 1156 675 1172
rect 641 164 675 180
rect 741 1138 821 1168
rect 741 198 761 1138
rect 801 300 821 1138
rect 801 200 1074 300
rect 801 198 821 200
rect 741 168 821 198
rect -607 94 -51 114
rect -607 34 -587 94
rect -71 34 -51 94
rect -607 14 -51 34
rect 51 -34 607 -14
rect 51 -94 71 -34
rect 587 -94 607 -34
rect 51 -114 607 -94
rect -1074 -1318 -1054 -200
rect -1014 -1318 -994 -200
rect -841 -198 -761 -168
rect -841 -1138 -821 -198
rect -781 -1138 -761 -198
rect -841 -1168 -761 -1138
rect -675 -180 -641 -164
rect -675 -1172 -641 -1156
rect -17 -180 17 -164
rect -17 -1172 17 -1156
rect 641 -180 675 -164
rect 641 -1172 675 -1156
rect 761 -198 841 -168
rect 761 -1138 781 -198
rect 821 -1138 841 -198
rect 761 -1168 841 -1138
rect 994 -200 1074 200
rect -1074 -1348 -994 -1318
rect -687 -1262 687 -1242
rect -687 -1302 -657 -1262
rect 657 -1302 687 -1262
rect -687 -1322 687 -1302
rect 994 -1318 1014 -200
rect 1054 -1318 1074 -200
rect 994 -1348 1074 -1318
rect -868 -1494 868 -1474
rect -868 -1534 -838 -1494
rect 838 -1534 868 -1494
rect -868 -1554 868 -1534
<< viali >>
rect -657 1242 657 1282
rect -801 198 -761 1138
rect -675 180 -641 1156
rect -17 180 17 1156
rect 641 180 675 1156
rect 761 198 801 1138
rect -587 34 -71 94
rect 71 -94 587 -34
rect -1054 -1318 -1014 -200
rect -821 -1138 -781 -198
rect -675 -1156 -641 -180
rect -17 -1156 17 -180
rect 641 -1156 675 -180
rect 781 -1138 821 -198
rect -657 -1302 657 -1262
rect 1014 -1318 1054 -200
rect -838 -1534 838 -1494
<< metal1 >>
rect -841 1282 841 1422
rect -841 1242 -657 1282
rect 657 1242 841 1282
rect -841 1222 841 1242
rect -841 1168 -681 1222
rect 681 1168 841 1222
rect -841 1156 -635 1168
rect -841 1138 -675 1156
rect -841 198 -801 1138
rect -761 198 -675 1138
rect -841 180 -675 198
rect -641 180 -635 1156
rect -841 168 -635 180
rect -23 1156 23 1168
rect -23 180 -17 1156
rect 17 180 23 1156
rect -23 114 23 180
rect 635 1156 841 1168
rect 635 180 641 1156
rect 675 1138 841 1156
rect 675 198 761 1138
rect 801 198 841 1138
rect 675 180 841 198
rect 635 168 841 180
rect -607 94 -51 114
rect -607 34 -587 94
rect -71 34 -51 94
rect -607 14 -51 34
rect -23 14 681 114
rect 51 -34 607 -14
rect 51 -94 71 -34
rect 587 -94 607 -34
rect 51 -114 607 -94
rect -1094 -200 -994 -170
rect -1094 -1318 -1054 -200
rect -1014 -1318 -994 -200
rect -1094 -1474 -994 -1318
rect -841 -180 -635 -168
rect -841 -198 -675 -180
rect -841 -1138 -821 -198
rect -781 -1138 -675 -198
rect -841 -1156 -675 -1138
rect -641 -1156 -635 -180
rect -841 -1168 -635 -1156
rect -23 -180 23 -168
rect -23 -1156 -17 -180
rect 17 -1156 23 -180
rect -23 -1168 23 -1156
rect 635 -180 681 14
rect 635 -1156 641 -180
rect 675 -1156 681 -180
rect 635 -1168 681 -1156
rect 761 -198 841 -168
rect 761 -1138 781 -198
rect 821 -1138 841 -198
rect -841 -1242 -681 -1168
rect 761 -1242 841 -1138
rect -841 -1262 841 -1242
rect -841 -1302 -657 -1262
rect 657 -1302 841 -1262
rect -841 -1342 841 -1302
rect 994 -200 1094 -170
rect 994 -1318 1014 -200
rect 1054 -1318 1094 -200
rect 994 -1474 1094 -1318
rect -1094 -1494 1094 -1474
rect -1094 -1534 -838 -1494
rect 838 -1534 1094 -1494
rect -1094 -1574 1094 -1534
<< labels >>
rlabel metal1 581 14 681 114 3 AND
rlabel metal1 -841 1322 -741 1422 1 VDD
rlabel metal1 51 -114 607 -14 3 A
rlabel metal1 -607 14 -51 114 7 B
rlabel metal1 -841 -1342 -741 -1242 5 GND
<< end >>
