magic
tech sky130A
magscale 1 2
timestamp 1700104495
<< checkpaint >>
rect -2312 4212 5632 4912
rect -2312 -3032 6852 4212
rect -1092 -3732 6852 -3032
<< nwell >>
rect 758 261 1834 915
<< pwell >>
rect 803 981 1762 1156
rect 3 38 3018 204
<< locali >>
rect 855 1100 913 1180
rect 760 920 994 961
rect 17 460 75 540
rect 251 215 574 263
rect 760 257 800 920
rect 1138 916 1268 962
rect 855 620 913 700
rect 855 460 913 540
rect 608 256 800 257
rect 2004 256 2284 262
rect 608 222 760 256
rect 794 222 800 256
rect 608 215 800 222
rect 2004 220 2172 256
rect 2206 220 2284 256
rect 2318 220 2598 262
rect 17 0 75 100
rect 855 0 913 100
rect 260 -114 340 -100
rect 260 -166 274 -114
rect 326 -166 340 -114
rect 260 -180 340 -166
rect 3520 -114 3600 -100
rect 3520 -166 3534 -114
rect 3586 -166 3600 -114
rect 3520 -180 3600 -166
rect 263 -560 305 -180
rect 3535 -560 3577 -180
<< viali >>
rect 166 215 200 249
rect 1458 922 1492 956
rect 1646 920 1680 960
rect 760 222 794 256
rect 1080 222 1114 256
rect 1694 220 1728 256
rect 1912 220 1946 256
rect 2172 220 2206 256
rect 2682 220 2716 256
rect 2866 220 2900 260
rect 274 -166 326 -114
rect 3534 -166 3586 -114
<< metal1 >>
rect 0 1128 3840 1224
rect 1406 988 1544 1008
rect 1406 890 1426 988
rect 1524 890 1544 988
rect 1620 960 1700 980
rect 1620 920 1646 960
rect 1680 920 1700 960
rect 1620 900 1700 920
rect 1406 870 1544 890
rect 0 660 3020 680
rect 0 520 150 660
rect 210 520 3020 660
rect 0 496 3020 520
rect 1090 358 2680 412
rect 0 249 220 280
rect 1090 276 1136 358
rect 2630 308 2676 358
rect 0 215 166 249
rect 200 215 220 249
rect 0 200 220 215
rect 740 256 1136 276
rect 740 222 760 256
rect 794 222 1080 256
rect 1114 222 1136 256
rect 740 202 1136 222
rect 1090 198 1136 202
rect 1642 288 1780 308
rect 1642 188 1662 288
rect 1760 188 1780 288
rect 1642 170 1780 188
rect 1860 288 1998 308
rect 1860 188 1880 288
rect 1978 188 1998 288
rect 1860 170 1998 188
rect 2120 288 2258 308
rect 2120 188 2140 288
rect 2238 188 2258 288
rect 2120 170 2258 188
rect 2630 256 2768 308
rect 2630 220 2682 256
rect 2716 220 2768 256
rect 2630 170 2768 220
rect 2840 260 2920 280
rect 2840 220 2866 260
rect 2900 220 2920 260
rect 2840 200 2920 220
rect 0 -48 3020 48
rect 3740 -60 3840 1128
rect 260 -114 340 -100
rect 260 -166 274 -114
rect 326 -166 340 -114
rect 260 -180 340 -166
rect 3520 -114 3600 -100
rect 3520 -166 3534 -114
rect 3586 -166 3600 -114
rect 3520 -180 3600 -166
<< via1 >>
rect 1426 956 1524 988
rect 1426 922 1458 956
rect 1458 922 1492 956
rect 1492 922 1524 956
rect 1426 890 1524 922
rect 150 520 210 660
rect 1662 256 1760 288
rect 1662 220 1694 256
rect 1694 220 1728 256
rect 1728 220 1760 256
rect 1662 188 1760 220
rect 1880 256 1978 288
rect 1880 220 1912 256
rect 1912 220 1946 256
rect 1946 220 1978 256
rect 1880 188 1978 220
rect 2140 256 2238 288
rect 2140 220 2172 256
rect 2172 220 2206 256
rect 2206 220 2238 256
rect 2140 188 2238 220
rect 274 -166 326 -114
rect 3534 -166 3586 -114
rect 564 -380 716 -320
rect 1844 -380 1996 -320
rect 3124 -380 3276 -320
<< metal2 >>
rect 1406 988 1544 1008
rect 1406 890 1426 988
rect 1524 890 1544 988
rect 1406 880 1544 890
rect 1406 870 2208 880
rect 1421 840 2208 870
rect 130 660 230 680
rect 130 520 150 660
rect 210 520 230 660
rect 130 -300 230 520
rect 2172 308 2208 840
rect 1642 288 1780 308
rect 1642 188 1662 288
rect 1760 188 1780 288
rect 1642 170 1780 188
rect 1860 288 1998 308
rect 1860 188 1880 288
rect 1978 188 1998 288
rect 1860 170 1998 188
rect 2120 288 2258 308
rect 2120 188 2140 288
rect 2238 188 2258 288
rect 2120 170 2258 188
rect 1680 -100 1740 170
rect 260 -114 1740 -100
rect 260 -166 274 -114
rect 326 -160 1740 -114
rect 1900 -100 1960 170
rect 1900 -114 3600 -100
rect 1900 -160 3534 -114
rect 326 -166 340 -160
rect 260 -180 340 -166
rect 3520 -166 3534 -160
rect 3586 -166 3600 -114
rect 3520 -180 3600 -166
rect 130 -320 3300 -300
rect 130 -380 564 -320
rect 716 -380 1844 -320
rect 1996 -380 3124 -320
rect 3276 -380 3300 -320
rect 130 -400 3300 -380
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2468 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_1
timestamp 1683767628
transform 1 0 1244 0 -1 1176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 444 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1683767628
transform 1 0 1840 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1683767628
transform 1 0 2154 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1683767628
transform 1 0 930 0 -1 1176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 130 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 930 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 0 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_1
timestamp 1683767628
transform 1 0 838 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_2
timestamp 1683767628
transform 1 0 838 0 -1 1176
box -38 -48 130 592
use sp_delay_top  sp_delay_top_0
timestamp 1700082107
transform 0 1 0 -1 0 42
box 0 0 6422 3840
<< labels >>
rlabel metal1 3740 1100 3840 1200 1 VSS
port 1 n
rlabel metal2 130 580 230 680 1 VCC
port 2 n
rlabel metal1 0 200 80 280 7 Vin
port 3 w
rlabel metal1 1620 900 1700 980 3 VFE
port 4 e
rlabel metal1 2840 200 2920 280 3 VRE
port 5 e
<< end >>
