magic
tech sky130A
magscale 1 2
timestamp 1699934371
<< dnwell >>
rect -187 -1532 7721 108
<< nwell >>
rect -267 -98 7801 2502
rect -267 -1326 19 -98
rect 7515 -1326 7801 -98
rect -267 -1612 7801 -1326
<< pwell >>
rect 19 -1326 7515 -98
<< mvnsubdiff >>
rect -187 -196 -107 -166
rect -187 -1296 -167 -196
rect -127 -1296 -107 -196
rect -187 -1326 -107 -1296
rect 7641 -196 7721 -166
rect 7641 -1296 7661 -196
rect 7701 -1296 7721 -196
rect 7641 -1326 7721 -1296
rect 19 -1472 7515 -1452
rect 19 -1512 49 -1472
rect 7485 -1512 7515 -1472
rect 19 -1532 7515 -1512
<< mvnsubdiffcont >>
rect -167 -1296 -127 -196
rect 7661 -1296 7701 -196
rect 49 -1512 7485 -1472
<< locali >>
rect -187 200 99 300
rect 7435 200 7721 300
rect -187 -196 -107 200
rect -187 -1296 -167 -196
rect -127 -1296 -107 -196
rect -187 -1326 -107 -1296
rect 7641 -196 7721 200
rect 7641 -1296 7661 -196
rect 7701 -1296 7721 -196
rect 7641 -1326 7721 -1296
rect 19 -1472 7515 -1452
rect 19 -1512 49 -1472
rect 7485 -1512 7515 -1472
rect 19 -1532 7515 -1512
<< viali >>
rect -167 -1296 -127 -196
rect 7661 -1296 7701 -196
rect 49 -1512 7485 -1472
<< metal1 >>
rect -3586 2400 7468 2600
rect 660 1460 1060 2400
rect 2500 1460 2900 2400
rect 66 1260 4340 1460
rect 1400 16 2200 116
rect 3200 96 3680 116
rect 3296 36 3680 96
rect 3200 16 3680 36
rect -834 -32 1140 -12
rect -834 -92 -814 -32
rect -754 -92 1140 -32
rect -834 -112 1140 -92
rect -207 -196 -107 -166
rect -207 -1296 -167 -196
rect -127 -1296 -107 -196
rect 1738 -1060 1838 16
rect 3580 -824 3680 16
rect 3580 -884 3600 -824
rect 3660 -884 3680 -824
rect 3580 -904 3680 -884
rect 7641 -196 7741 -166
rect 1738 -1120 1758 -1060
rect 1818 -1120 1838 -1060
rect 1738 -1140 1838 -1120
rect 3730 -1076 4320 -980
rect 3730 -1220 7488 -1076
rect -207 -1452 -107 -1296
rect 46 -1300 7488 -1220
rect 7641 -1296 7661 -196
rect 7701 -1296 7741 -196
rect 7641 -1452 7741 -1296
rect -542 -1472 7741 -1452
rect -542 -1512 49 -1472
rect 7485 -1512 7741 -1472
rect -542 -1552 7741 -1512
rect -542 -1652 7408 -1552
<< via1 >>
rect 280 36 796 96
rect 2780 36 3296 96
rect -814 -92 -754 -32
rect 2780 -92 3296 -32
rect 3600 -884 3660 -824
rect 1758 -1120 1818 -1060
<< metal2 >>
rect -1734 1118 -594 1218
rect -1734 990 -734 1090
rect -834 -32 -734 990
rect -834 -92 -814 -32
rect -754 -92 -734 -32
rect -834 -112 -734 -92
rect -694 -12 -594 1118
rect 260 96 3316 116
rect 260 36 280 96
rect 796 36 2780 96
rect 3296 36 3316 96
rect 260 16 3316 36
rect -694 -32 3316 -12
rect -694 -92 2780 -32
rect 3296 -92 3316 -32
rect -694 -112 3316 -92
rect 3580 -824 4000 -804
rect 3580 -884 3600 -824
rect 3660 -884 4000 -824
rect 3580 -904 4000 -884
rect 1738 -1060 1838 -1040
rect 1738 -1120 1758 -1060
rect 1818 -1120 1838 -1060
rect 1738 -1300 1838 -1120
rect 4102 -1300 4202 -804
rect 1738 -1400 4202 -1300
use boot_ls_stage  boot_ls_stage_0
timestamp 1699931927
transform 1 0 -2811 0 1 1104
box -1778 -2264 1444 1422
use buffer  buffer_0
timestamp 1699046184
transform 1 0 4051 0 1 -12
box -395 -1088 3503 2502
use nand_5v  nand_5v_0
timestamp 1699045454
transform 1 0 867 0 1 2
box -867 -1302 867 1348
use nand_5v  nand_5v_1
timestamp 1699045454
transform 1 0 2709 0 1 2
box -867 -1302 867 1348
<< labels >>
rlabel metal1 -3586 2400 -3386 2600 1 VBOOT
rlabel metal1 7208 -1652 7408 -1452 5 VSource
<< end >>
