magic
tech sky130A
magscale 1 2
timestamp 1699035782
<< dnwell >>
rect -554 -1214 3704 120
rect 28 -1340 3704 -1214
<< nwell >>
rect 215 954 3517 2522
rect -395 200 3517 954
rect -634 -86 3784 200
rect -634 -1008 -348 -86
rect -634 -1134 234 -1008
rect 3498 -1134 3784 -86
rect -634 -1294 3784 -1134
rect -52 -1420 3784 -1294
<< pwell >>
rect -348 -1008 3498 -86
rect 234 -1134 3498 -1008
<< mvnmos >>
rect -129 -754 -29 -154
rect 29 -754 129 -154
rect 473 -954 573 -154
rect 631 -954 731 -154
rect 789 -954 889 -154
rect 947 -954 1047 -154
rect 1105 -954 1205 -154
rect 1263 -954 1363 -154
rect 1421 -954 1521 -154
rect 1579 -954 1679 -154
rect 1737 -954 1837 -154
rect 1895 -954 1995 -154
rect 2053 -954 2153 -154
rect 2211 -954 2311 -154
rect 2369 -954 2469 -154
rect 2527 -954 2627 -154
rect 2685 -954 2785 -154
rect 2843 -954 2943 -154
rect 3001 -954 3101 -154
rect 3159 -954 3259 -154
<< mvpmos >>
rect -137 154 -37 354
rect 37 154 137 754
rect 473 154 573 2322
rect 631 154 731 2322
rect 789 154 889 2322
rect 947 154 1047 2322
rect 1105 154 1205 2322
rect 1263 154 1363 2322
rect 1421 154 1521 2322
rect 1579 154 1679 2322
rect 1737 154 1837 2322
rect 1895 154 1995 2322
rect 2053 154 2153 2322
rect 2211 154 2311 2322
rect 2369 154 2469 2322
rect 2527 154 2627 2322
rect 2685 154 2785 2322
rect 2843 154 2943 2322
rect 3001 154 3101 2322
rect 3159 154 3259 2322
<< mvndiff >>
rect -187 -166 -129 -154
rect -187 -742 -175 -166
rect -141 -742 -129 -166
rect -187 -754 -129 -742
rect -29 -166 29 -154
rect -29 -742 -17 -166
rect 17 -742 29 -166
rect -29 -754 29 -742
rect 129 -166 187 -154
rect 129 -742 141 -166
rect 175 -742 187 -166
rect 129 -754 187 -742
rect 415 -166 473 -154
rect 415 -942 427 -166
rect 461 -942 473 -166
rect 415 -954 473 -942
rect 573 -166 631 -154
rect 573 -942 585 -166
rect 619 -942 631 -166
rect 573 -954 631 -942
rect 731 -166 789 -154
rect 731 -942 743 -166
rect 777 -942 789 -166
rect 731 -954 789 -942
rect 889 -166 947 -154
rect 889 -942 901 -166
rect 935 -942 947 -166
rect 889 -954 947 -942
rect 1047 -166 1105 -154
rect 1047 -942 1059 -166
rect 1093 -942 1105 -166
rect 1047 -954 1105 -942
rect 1205 -166 1263 -154
rect 1205 -942 1217 -166
rect 1251 -942 1263 -166
rect 1205 -954 1263 -942
rect 1363 -166 1421 -154
rect 1363 -942 1375 -166
rect 1409 -942 1421 -166
rect 1363 -954 1421 -942
rect 1521 -166 1579 -154
rect 1521 -942 1533 -166
rect 1567 -942 1579 -166
rect 1521 -954 1579 -942
rect 1679 -166 1737 -154
rect 1679 -942 1691 -166
rect 1725 -942 1737 -166
rect 1679 -954 1737 -942
rect 1837 -166 1895 -154
rect 1837 -942 1849 -166
rect 1883 -942 1895 -166
rect 1837 -954 1895 -942
rect 1995 -166 2053 -154
rect 1995 -942 2007 -166
rect 2041 -942 2053 -166
rect 1995 -954 2053 -942
rect 2153 -166 2211 -154
rect 2153 -942 2165 -166
rect 2199 -942 2211 -166
rect 2153 -954 2211 -942
rect 2311 -166 2369 -154
rect 2311 -942 2323 -166
rect 2357 -942 2369 -166
rect 2311 -954 2369 -942
rect 2469 -166 2527 -154
rect 2469 -942 2481 -166
rect 2515 -942 2527 -166
rect 2469 -954 2527 -942
rect 2627 -166 2685 -154
rect 2627 -942 2639 -166
rect 2673 -942 2685 -166
rect 2627 -954 2685 -942
rect 2785 -166 2843 -154
rect 2785 -942 2797 -166
rect 2831 -942 2843 -166
rect 2785 -954 2843 -942
rect 2943 -166 3001 -154
rect 2943 -942 2955 -166
rect 2989 -942 3001 -166
rect 2943 -954 3001 -942
rect 3101 -166 3159 -154
rect 3101 -942 3113 -166
rect 3147 -942 3159 -166
rect 3101 -954 3159 -942
rect 3259 -166 3317 -154
rect 3259 -942 3271 -166
rect 3305 -942 3317 -166
rect 3259 -954 3317 -942
<< mvpdiff >>
rect -21 742 37 754
rect -21 354 -9 742
rect -195 342 -137 354
rect -195 166 -183 342
rect -149 166 -137 342
rect -195 154 -137 166
rect -37 342 -9 354
rect -37 166 -25 342
rect 25 166 37 742
rect -37 154 37 166
rect 137 742 195 754
rect 137 166 149 742
rect 183 166 195 742
rect 137 154 195 166
rect 415 2310 473 2322
rect 415 166 427 2310
rect 461 166 473 2310
rect 415 154 473 166
rect 573 2310 631 2322
rect 573 166 585 2310
rect 619 166 631 2310
rect 573 154 631 166
rect 731 2310 789 2322
rect 731 166 743 2310
rect 777 166 789 2310
rect 731 154 789 166
rect 889 2310 947 2322
rect 889 166 901 2310
rect 935 166 947 2310
rect 889 154 947 166
rect 1047 2310 1105 2322
rect 1047 166 1059 2310
rect 1093 166 1105 2310
rect 1047 154 1105 166
rect 1205 2310 1263 2322
rect 1205 166 1217 2310
rect 1251 166 1263 2310
rect 1205 154 1263 166
rect 1363 2310 1421 2322
rect 1363 166 1375 2310
rect 1409 166 1421 2310
rect 1363 154 1421 166
rect 1521 2310 1579 2322
rect 1521 166 1533 2310
rect 1567 166 1579 2310
rect 1521 154 1579 166
rect 1679 2310 1737 2322
rect 1679 166 1691 2310
rect 1725 166 1737 2310
rect 1679 154 1737 166
rect 1837 2310 1895 2322
rect 1837 166 1849 2310
rect 1883 166 1895 2310
rect 1837 154 1895 166
rect 1995 2310 2053 2322
rect 1995 166 2007 2310
rect 2041 166 2053 2310
rect 1995 154 2053 166
rect 2153 2310 2211 2322
rect 2153 166 2165 2310
rect 2199 166 2211 2310
rect 2153 154 2211 166
rect 2311 2310 2369 2322
rect 2311 166 2323 2310
rect 2357 166 2369 2310
rect 2311 154 2369 166
rect 2469 2310 2527 2322
rect 2469 166 2481 2310
rect 2515 166 2527 2310
rect 2469 154 2527 166
rect 2627 2310 2685 2322
rect 2627 166 2639 2310
rect 2673 166 2685 2310
rect 2627 154 2685 166
rect 2785 2310 2843 2322
rect 2785 166 2797 2310
rect 2831 166 2843 2310
rect 2785 154 2843 166
rect 2943 2310 3001 2322
rect 2943 166 2955 2310
rect 2989 166 3001 2310
rect 2943 154 3001 166
rect 3101 2310 3159 2322
rect 3101 166 3113 2310
rect 3147 166 3159 2310
rect 3101 154 3159 166
rect 3259 2310 3317 2322
rect 3259 166 3271 2310
rect 3305 166 3317 2310
rect 3259 154 3317 166
<< mvndiffc >>
rect -175 -742 -141 -166
rect -17 -742 17 -166
rect 141 -742 175 -166
rect 427 -942 461 -166
rect 585 -942 619 -166
rect 743 -942 777 -166
rect 901 -942 935 -166
rect 1059 -942 1093 -166
rect 1217 -942 1251 -166
rect 1375 -942 1409 -166
rect 1533 -942 1567 -166
rect 1691 -942 1725 -166
rect 1849 -942 1883 -166
rect 2007 -942 2041 -166
rect 2165 -942 2199 -166
rect 2323 -942 2357 -166
rect 2481 -942 2515 -166
rect 2639 -942 2673 -166
rect 2797 -942 2831 -166
rect 2955 -942 2989 -166
rect 3113 -942 3147 -166
rect 3271 -942 3305 -166
<< mvpdiffc >>
rect -183 166 -149 342
rect -9 342 25 742
rect -25 166 25 342
rect 149 166 183 742
rect 427 166 461 2310
rect 585 166 619 2310
rect 743 166 777 2310
rect 901 166 935 2310
rect 1059 166 1093 2310
rect 1217 166 1251 2310
rect 1375 166 1409 2310
rect 1533 166 1567 2310
rect 1691 166 1725 2310
rect 1849 166 1883 2310
rect 2007 166 2041 2310
rect 2165 166 2199 2310
rect 2323 166 2357 2310
rect 2481 166 2515 2310
rect 2639 166 2673 2310
rect 2797 166 2831 2310
rect 2955 166 2989 2310
rect 3113 166 3147 2310
rect 3271 166 3305 2310
<< mvpsubdiff >>
rect -301 -184 -261 -154
rect -301 -754 -261 -724
rect 261 -184 341 -154
rect 261 -924 281 -184
rect 321 -924 341 -184
rect -187 -982 -157 -942
rect 157 -982 187 -942
rect 261 -954 341 -924
rect 3391 -184 3471 -154
rect 3391 -924 3411 -184
rect 3451 -924 3471 -184
rect 3391 -954 3471 -924
rect 415 -1048 3317 -1028
rect 415 -1088 445 -1048
rect 3287 -1088 3317 -1048
rect 415 -1108 3317 -1088
<< mvnsubdiff >>
rect 415 2436 3317 2456
rect 415 2396 445 2436
rect 3287 2396 3317 2436
rect 415 2376 3317 2396
rect 281 2292 361 2322
rect -195 808 -165 848
rect 165 808 195 848
rect -289 724 -249 754
rect -289 154 -249 184
rect 281 184 301 2292
rect 341 184 361 2292
rect 281 154 361 184
rect 3371 2292 3451 2322
rect 3371 184 3391 2292
rect 3431 184 3451 2292
rect 3371 154 3451 184
rect -514 -186 -474 -156
rect -514 -1008 -474 -978
rect 3624 -186 3704 -156
rect 3624 -1104 3644 -186
rect 3684 -1104 3704 -186
rect 3624 -1134 3704 -1104
rect -348 -1174 -318 -1134
rect 138 -1174 168 -1134
rect 234 -1280 3498 -1260
rect 234 -1320 264 -1280
rect 3468 -1320 3498 -1280
rect 234 -1340 3498 -1320
<< mvpsubdiffcont >>
rect -301 -724 -261 -184
rect 281 -924 321 -184
rect -157 -982 157 -942
rect 3411 -924 3451 -184
rect 445 -1088 3287 -1048
<< mvnsubdiffcont >>
rect 445 2396 3287 2436
rect -165 808 165 848
rect -289 184 -249 724
rect 301 184 341 2292
rect 3391 184 3431 2292
rect -514 -978 -474 -186
rect 3644 -1104 3684 -186
rect -318 -1174 138 -1134
rect 264 -1320 3468 -1280
<< poly >>
rect 473 2322 573 2348
rect 631 2322 731 2348
rect 789 2322 889 2348
rect 947 2322 1047 2348
rect 1105 2322 1205 2348
rect 1263 2322 1363 2348
rect 1421 2322 1521 2348
rect 1579 2322 1679 2348
rect 1737 2322 1837 2348
rect 1895 2322 1995 2348
rect 2053 2322 2153 2348
rect 2211 2322 2311 2348
rect 2369 2322 2469 2348
rect 2527 2322 2627 2348
rect 2685 2322 2785 2348
rect 2843 2322 2943 2348
rect 3001 2322 3101 2348
rect 3159 2322 3259 2348
rect 37 754 137 780
rect -137 354 -37 380
rect -137 96 -37 154
rect -137 36 -117 96
rect -57 36 -37 96
rect -137 16 -37 36
rect 37 96 137 154
rect 37 36 57 96
rect 117 36 137 96
rect 37 16 137 36
rect 473 -14 573 154
rect 449 -34 573 -14
rect 449 -94 469 -34
rect 529 -94 573 -34
rect 449 -114 573 -94
rect -129 -154 -29 -128
rect 29 -154 129 -128
rect 473 -154 573 -114
rect 631 -14 731 154
rect 789 -14 889 154
rect 631 -34 889 -14
rect 631 -94 675 -34
rect 845 -94 889 -34
rect 631 -114 889 -94
rect 631 -154 731 -114
rect 789 -154 889 -114
rect 947 -14 1047 154
rect 1105 -14 1205 154
rect 947 -34 1205 -14
rect 947 -94 991 -34
rect 1161 -94 1205 -34
rect 947 -114 1205 -94
rect 947 -154 1047 -114
rect 1105 -154 1205 -114
rect 1263 -14 1363 154
rect 1421 -14 1521 154
rect 1263 -34 1521 -14
rect 1263 -94 1307 -34
rect 1477 -94 1521 -34
rect 1263 -114 1521 -94
rect 1263 -154 1363 -114
rect 1421 -154 1521 -114
rect 1579 -14 1679 154
rect 1737 -14 1837 154
rect 1579 -34 1837 -14
rect 1579 -94 1623 -34
rect 1793 -94 1837 -34
rect 1579 -114 1837 -94
rect 1579 -154 1679 -114
rect 1737 -154 1837 -114
rect 1895 -14 1995 154
rect 2053 -14 2153 154
rect 1895 -34 2153 -14
rect 1895 -94 1939 -34
rect 2109 -94 2153 -34
rect 1895 -114 2153 -94
rect 1895 -154 1995 -114
rect 2053 -154 2153 -114
rect 2211 -14 2311 154
rect 2369 -14 2469 154
rect 2211 -34 2469 -14
rect 2211 -94 2255 -34
rect 2425 -94 2469 -34
rect 2211 -114 2469 -94
rect 2211 -154 2311 -114
rect 2369 -154 2469 -114
rect 2527 -14 2627 154
rect 2685 -14 2785 154
rect 2527 -34 2785 -14
rect 2527 -94 2571 -34
rect 2741 -94 2785 -34
rect 2527 -114 2785 -94
rect 2527 -154 2627 -114
rect 2685 -154 2785 -114
rect 2843 -14 2943 154
rect 3001 -14 3101 154
rect 2843 -34 3101 -14
rect 2843 -94 2887 -34
rect 3057 -94 3101 -34
rect 2843 -114 3101 -94
rect 2843 -154 2943 -114
rect 3001 -154 3101 -114
rect 3159 -14 3259 154
rect 3159 -34 3283 -14
rect 3159 -94 3203 -34
rect 3263 -94 3283 -34
rect 3159 -114 3283 -94
rect 3159 -154 3259 -114
rect -129 -812 -29 -754
rect -129 -872 -109 -812
rect -49 -872 -29 -812
rect -129 -892 -29 -872
rect 29 -812 129 -754
rect 29 -872 49 -812
rect 109 -872 129 -812
rect 29 -892 129 -872
rect 473 -980 573 -954
rect 631 -980 731 -954
rect 789 -980 889 -954
rect 947 -980 1047 -954
rect 1105 -980 1205 -954
rect 1263 -980 1363 -954
rect 1421 -980 1521 -954
rect 1579 -980 1679 -954
rect 1737 -980 1837 -954
rect 1895 -980 1995 -954
rect 2053 -980 2153 -954
rect 2211 -980 2311 -954
rect 2369 -980 2469 -954
rect 2527 -980 2627 -954
rect 2685 -980 2785 -954
rect 2843 -980 2943 -954
rect 3001 -980 3101 -954
rect 3159 -980 3259 -954
<< polycont >>
rect -117 36 -57 96
rect 57 36 117 96
rect 469 -94 529 -34
rect 675 -94 845 -34
rect 991 -94 1161 -34
rect 1307 -94 1477 -34
rect 1623 -94 1793 -34
rect 1939 -94 2109 -34
rect 2255 -94 2425 -34
rect 2571 -94 2741 -34
rect 2887 -94 3057 -34
rect 3203 -94 3263 -34
rect -109 -872 -49 -812
rect 49 -872 109 -812
<< locali >>
rect 415 2436 3317 2456
rect 415 2396 445 2436
rect 3287 2396 3317 2436
rect 415 2376 3317 2396
rect 281 2292 361 2322
rect -195 808 -165 848
rect 165 808 195 848
rect -289 724 -249 754
rect -9 742 25 758
rect -289 154 -249 184
rect -183 342 -149 358
rect -183 150 -149 166
rect -25 342 -9 358
rect -25 150 25 166
rect 149 742 183 758
rect 149 150 183 166
rect 281 184 301 2292
rect 341 184 361 2292
rect 281 154 361 184
rect 427 2310 461 2326
rect 427 150 461 166
rect 585 2310 619 2326
rect 585 150 619 166
rect 743 2310 777 2326
rect 743 150 777 166
rect 901 2310 935 2326
rect 901 150 935 166
rect 1059 2310 1093 2326
rect 1059 150 1093 166
rect 1217 2310 1251 2326
rect 1217 150 1251 166
rect 1375 2310 1409 2326
rect 1375 150 1409 166
rect 1533 2310 1567 2326
rect 1533 150 1567 166
rect 1691 2310 1725 2326
rect 1691 150 1725 166
rect 1849 2310 1883 2326
rect 1849 150 1883 166
rect 2007 2310 2041 2326
rect 2007 150 2041 166
rect 2165 2310 2199 2326
rect 2165 150 2199 166
rect 2323 2310 2357 2326
rect 2323 150 2357 166
rect 2481 2310 2515 2326
rect 2481 150 2515 166
rect 2639 2310 2673 2326
rect 2639 150 2673 166
rect 2797 2310 2831 2326
rect 2797 150 2831 166
rect 2955 2310 2989 2326
rect 2955 150 2989 166
rect 3113 2310 3147 2326
rect 3113 150 3147 166
rect 3271 2310 3305 2326
rect 3271 150 3305 166
rect 3371 2292 3451 2322
rect 3371 184 3391 2292
rect 3431 254 3451 2292
rect 3431 184 3704 254
rect 3371 154 3704 184
rect -137 96 -37 116
rect -137 36 -117 96
rect -57 36 -37 96
rect -137 -16 -37 36
rect 7 96 137 116
rect 7 36 27 96
rect 117 36 137 96
rect 7 16 137 36
rect -137 -36 -7 -16
rect -137 -96 -87 -36
rect -27 -96 -7 -36
rect -137 -116 -7 -96
rect 449 -34 549 -14
rect 449 -94 469 -34
rect 529 -94 549 -34
rect 449 -114 549 -94
rect 655 -34 865 -14
rect 655 -94 675 -34
rect 845 -94 865 -34
rect 655 -114 865 -94
rect 971 -34 1181 -14
rect 971 -94 991 -34
rect 1161 -94 1181 -34
rect 971 -114 1181 -94
rect 1287 -34 1497 -14
rect 1287 -94 1307 -34
rect 1477 -94 1497 -34
rect 1287 -114 1497 -94
rect 1603 -34 1813 -14
rect 1603 -94 1623 -34
rect 1793 -94 1813 -34
rect 1603 -114 1813 -94
rect 1919 -34 2129 -14
rect 1919 -94 1939 -34
rect 2109 -94 2129 -34
rect 1919 -114 2129 -94
rect 2235 -34 2445 -14
rect 2235 -94 2255 -34
rect 2425 -94 2445 -34
rect 2235 -114 2445 -94
rect 2551 -34 2761 -14
rect 2551 -94 2571 -34
rect 2741 -94 2761 -34
rect 2551 -114 2761 -94
rect 2867 -34 3077 -14
rect 2867 -94 2887 -34
rect 3057 -94 3077 -34
rect 2867 -114 3077 -94
rect 3183 -34 3283 -14
rect 3183 -94 3203 -34
rect 3263 -94 3283 -34
rect 3183 -114 3283 -94
rect -514 -186 -474 -156
rect -301 -184 -261 -154
rect -301 -754 -261 -724
rect -175 -166 -141 -150
rect -175 -758 -141 -742
rect -17 -166 17 -150
rect -17 -758 17 -742
rect 141 -166 175 -150
rect 141 -758 175 -742
rect 261 -184 341 -154
rect -151 -812 -29 -792
rect -151 -872 -131 -812
rect -49 -872 -29 -812
rect -151 -892 -29 -872
rect 29 -812 151 -792
rect 29 -872 49 -812
rect 131 -872 151 -812
rect 29 -892 151 -872
rect 261 -924 281 -184
rect 321 -924 341 -184
rect -514 -1008 -474 -978
rect -187 -982 -157 -942
rect 157 -982 187 -942
rect 261 -954 341 -924
rect 427 -166 461 -150
rect 427 -958 461 -942
rect 585 -166 619 -150
rect 585 -958 619 -942
rect 743 -166 777 -150
rect 743 -958 777 -942
rect 901 -166 935 -150
rect 901 -958 935 -942
rect 1059 -166 1093 -150
rect 1059 -958 1093 -942
rect 1217 -166 1251 -150
rect 1217 -958 1251 -942
rect 1375 -166 1409 -150
rect 1375 -958 1409 -942
rect 1533 -166 1567 -150
rect 1533 -958 1567 -942
rect 1691 -166 1725 -150
rect 1691 -958 1725 -942
rect 1849 -166 1883 -150
rect 1849 -958 1883 -942
rect 2007 -166 2041 -150
rect 2007 -958 2041 -942
rect 2165 -166 2199 -150
rect 2165 -958 2199 -942
rect 2323 -166 2357 -150
rect 2323 -958 2357 -942
rect 2481 -166 2515 -150
rect 2481 -958 2515 -942
rect 2639 -166 2673 -150
rect 2639 -958 2673 -942
rect 2797 -166 2831 -150
rect 2797 -958 2831 -942
rect 2955 -166 2989 -150
rect 2955 -958 2989 -942
rect 3113 -166 3147 -150
rect 3113 -958 3147 -942
rect 3271 -166 3305 -150
rect 3271 -958 3305 -942
rect 3391 -184 3471 -154
rect 3391 -924 3411 -184
rect 3451 -924 3471 -184
rect 3391 -954 3471 -924
rect 3624 -186 3704 154
rect 415 -1048 3317 -1028
rect 415 -1088 445 -1048
rect 3287 -1088 3317 -1048
rect 415 -1108 3317 -1088
rect 3624 -1104 3644 -186
rect 3684 -1104 3704 -186
rect 3624 -1134 3704 -1104
rect -348 -1174 -318 -1134
rect 138 -1174 168 -1134
rect 234 -1280 3498 -1260
rect 234 -1320 264 -1280
rect 3468 -1320 3498 -1280
rect 234 -1340 3498 -1320
<< viali >>
rect 445 2396 3287 2436
rect -165 808 165 848
rect -289 184 -249 724
rect -183 166 -149 342
rect -9 342 25 742
rect -25 166 25 342
rect 149 166 183 742
rect 301 184 341 2292
rect 427 166 461 2310
rect 585 166 619 2310
rect 743 166 777 2310
rect 901 166 935 2310
rect 1059 166 1093 2310
rect 1217 166 1251 2310
rect 1375 166 1409 2310
rect 1533 166 1567 2310
rect 1691 166 1725 2310
rect 1849 166 1883 2310
rect 2007 166 2041 2310
rect 2165 166 2199 2310
rect 2323 166 2357 2310
rect 2481 166 2515 2310
rect 2639 166 2673 2310
rect 2797 166 2831 2310
rect 2955 166 2989 2310
rect 3113 166 3147 2310
rect 3271 166 3305 2310
rect 3391 184 3431 2292
rect 27 36 57 96
rect 57 36 87 96
rect -87 -96 -27 -36
rect 469 -94 529 -34
rect 675 -94 845 -34
rect 991 -94 1161 -34
rect 1307 -94 1477 -34
rect 1623 -94 1793 -34
rect 1939 -94 2109 -34
rect 2255 -94 2425 -34
rect 2571 -94 2741 -34
rect 2887 -94 3057 -34
rect 3203 -94 3263 -34
rect -514 -978 -474 -186
rect -301 -724 -261 -184
rect -175 -742 -141 -166
rect -17 -742 17 -166
rect 141 -742 175 -166
rect -131 -872 -109 -812
rect -109 -872 -71 -812
rect 71 -872 109 -812
rect 109 -872 131 -812
rect 281 -924 321 -184
rect -157 -982 157 -942
rect 427 -942 461 -166
rect 585 -942 619 -166
rect 743 -942 777 -166
rect 901 -942 935 -166
rect 1059 -942 1093 -166
rect 1217 -942 1251 -166
rect 1375 -942 1409 -166
rect 1533 -942 1567 -166
rect 1691 -942 1725 -166
rect 1849 -942 1883 -166
rect 2007 -942 2041 -166
rect 2165 -942 2199 -166
rect 2323 -942 2357 -166
rect 2481 -942 2515 -166
rect 2639 -942 2673 -166
rect 2797 -942 2831 -166
rect 2955 -942 2989 -166
rect 3113 -942 3147 -166
rect 3271 -942 3305 -166
rect 3411 -924 3451 -184
rect 445 -1088 3287 -1048
rect 3644 -1104 3684 -186
rect -318 -1174 138 -1134
rect 264 -1320 3468 -1280
<< metal1 >>
rect 261 2436 3471 2576
rect 261 2396 445 2436
rect 3287 2396 3471 2436
rect 261 2376 3471 2396
rect 261 2310 467 2376
rect 261 2292 427 2310
rect 261 988 301 2292
rect -309 848 301 988
rect -309 808 -165 848
rect 165 808 301 848
rect -309 788 301 808
rect -309 724 -229 788
rect -309 300 -289 724
rect -554 200 -289 300
rect -554 -186 -454 200
rect -309 184 -289 200
rect -249 184 -229 724
rect -15 742 31 788
rect -15 354 -9 742
rect -309 154 -229 184
rect -189 342 -143 354
rect -189 166 -183 342
rect -149 166 -143 342
rect -189 116 -143 166
rect -31 342 -9 354
rect -31 166 -25 342
rect 25 166 31 742
rect -31 154 31 166
rect 143 742 189 754
rect 143 166 149 742
rect 183 166 189 742
rect -189 96 107 116
rect -189 36 27 96
rect 87 36 107 96
rect -189 16 107 36
rect -554 -978 -514 -186
rect -474 -978 -454 -186
rect -554 -1114 -454 -978
rect -321 -184 -241 -154
rect -321 -724 -301 -184
rect -261 -724 -241 -184
rect -321 -922 -241 -724
rect -181 -166 -135 16
rect 143 -16 189 166
rect 261 184 301 788
rect 341 184 427 2292
rect 261 166 427 184
rect 461 166 467 2310
rect 261 154 467 166
rect 579 2310 625 2322
rect 579 166 585 2310
rect 619 166 625 2310
rect 579 114 625 166
rect 737 2310 783 2376
rect 737 166 743 2310
rect 777 166 783 2310
rect 737 154 783 166
rect 895 2310 941 2322
rect 895 166 901 2310
rect 935 166 941 2310
rect 895 114 941 166
rect 1053 2310 1099 2376
rect 1053 166 1059 2310
rect 1093 166 1099 2310
rect 1053 154 1099 166
rect 1211 2310 1257 2322
rect 1211 166 1217 2310
rect 1251 166 1257 2310
rect 1211 114 1257 166
rect 1369 2310 1415 2376
rect 1369 166 1375 2310
rect 1409 166 1415 2310
rect 1369 154 1415 166
rect 1527 2310 1573 2322
rect 1527 166 1533 2310
rect 1567 166 1573 2310
rect 1527 114 1573 166
rect 1685 2310 1731 2376
rect 1685 166 1691 2310
rect 1725 166 1731 2310
rect 1685 154 1731 166
rect 1843 2310 1889 2322
rect 1843 166 1849 2310
rect 1883 166 1889 2310
rect 1843 114 1889 166
rect 2001 2310 2047 2376
rect 2001 166 2007 2310
rect 2041 166 2047 2310
rect 2001 154 2047 166
rect 2159 2310 2205 2322
rect 2159 166 2165 2310
rect 2199 166 2205 2310
rect 2159 114 2205 166
rect 2317 2310 2363 2376
rect 2317 166 2323 2310
rect 2357 166 2363 2310
rect 2317 154 2363 166
rect 2475 2310 2521 2322
rect 2475 166 2481 2310
rect 2515 166 2521 2310
rect 2475 114 2521 166
rect 2633 2310 2679 2376
rect 2633 166 2639 2310
rect 2673 166 2679 2310
rect 2633 154 2679 166
rect 2791 2310 2837 2322
rect 2791 166 2797 2310
rect 2831 166 2837 2310
rect 2791 114 2837 166
rect 2949 2310 2995 2376
rect 2949 166 2955 2310
rect 2989 166 2995 2310
rect 2949 154 2995 166
rect 3107 2310 3153 2322
rect 3107 166 3113 2310
rect 3147 166 3153 2310
rect 3107 114 3153 166
rect 3265 2310 3471 2376
rect 3265 166 3271 2310
rect 3305 2292 3471 2310
rect 3305 184 3391 2292
rect 3431 184 3471 2292
rect 3305 166 3471 184
rect 3265 154 3471 166
rect 579 94 3153 114
rect 579 34 599 94
rect 3133 34 3153 94
rect 579 14 3153 34
rect -107 -36 189 -16
rect -107 -96 -87 -36
rect -27 -96 127 -36
rect 187 -96 189 -36
rect -107 -116 189 -96
rect 449 -34 549 -14
rect 449 -94 469 -34
rect 529 -94 549 -34
rect 449 -114 549 -94
rect -181 -742 -175 -166
rect -141 -742 -135 -166
rect -181 -754 -135 -742
rect -23 -166 23 -154
rect -23 -742 -17 -166
rect 17 -742 23 -166
rect -151 -812 -51 -792
rect -151 -872 -131 -812
rect -71 -872 -51 -812
rect -151 -892 -51 -872
rect -23 -922 23 -742
rect 135 -166 181 -116
rect 135 -742 141 -166
rect 175 -742 181 -166
rect 135 -754 181 -742
rect 261 -166 467 -154
rect 261 -184 427 -166
rect 51 -812 151 -792
rect 51 -872 71 -812
rect 131 -872 151 -812
rect 51 -892 151 -872
rect 261 -922 281 -184
rect -321 -924 281 -922
rect 321 -924 427 -184
rect -321 -942 427 -924
rect 461 -942 467 -166
rect -321 -982 -157 -942
rect 157 -982 467 -942
rect 579 -166 625 14
rect 655 -34 865 -14
rect 655 -94 675 -34
rect 845 -94 865 -34
rect 655 -114 865 -94
rect 579 -942 585 -166
rect 619 -942 625 -166
rect 579 -954 625 -942
rect 737 -166 783 -154
rect 737 -942 743 -166
rect 777 -942 783 -166
rect -321 -1002 467 -982
rect 261 -1028 467 -1002
rect 737 -1028 783 -942
rect 895 -166 941 14
rect 971 -34 1181 -14
rect 971 -94 991 -34
rect 1161 -94 1181 -34
rect 971 -114 1181 -94
rect 895 -942 901 -166
rect 935 -942 941 -166
rect 895 -954 941 -942
rect 1053 -166 1099 -154
rect 1053 -942 1059 -166
rect 1093 -942 1099 -166
rect 1053 -1028 1099 -942
rect 1211 -166 1257 14
rect 1287 -34 1497 -14
rect 1287 -94 1307 -34
rect 1477 -94 1497 -34
rect 1287 -114 1497 -94
rect 1211 -942 1217 -166
rect 1251 -942 1257 -166
rect 1211 -954 1257 -942
rect 1369 -166 1415 -154
rect 1369 -942 1375 -166
rect 1409 -942 1415 -166
rect 1369 -1028 1415 -942
rect 1527 -166 1573 14
rect 1603 -34 1813 -14
rect 1603 -94 1623 -34
rect 1793 -94 1813 -34
rect 1603 -114 1813 -94
rect 1527 -942 1533 -166
rect 1567 -942 1573 -166
rect 1527 -954 1573 -942
rect 1685 -166 1731 -154
rect 1685 -942 1691 -166
rect 1725 -942 1731 -166
rect 1685 -1028 1731 -942
rect 1843 -166 1889 14
rect 1919 -34 2129 -14
rect 1919 -94 1939 -34
rect 2109 -94 2129 -34
rect 1919 -114 2129 -94
rect 1843 -942 1849 -166
rect 1883 -942 1889 -166
rect 1843 -954 1889 -942
rect 2001 -166 2047 -154
rect 2001 -942 2007 -166
rect 2041 -942 2047 -166
rect 2001 -1028 2047 -942
rect 2159 -166 2205 14
rect 2235 -34 2445 -14
rect 2235 -94 2255 -34
rect 2425 -94 2445 -34
rect 2235 -114 2445 -94
rect 2159 -942 2165 -166
rect 2199 -942 2205 -166
rect 2159 -954 2205 -942
rect 2317 -166 2363 -154
rect 2317 -942 2323 -166
rect 2357 -942 2363 -166
rect 2317 -1028 2363 -942
rect 2475 -166 2521 14
rect 2551 -34 2761 -14
rect 2551 -94 2571 -34
rect 2741 -94 2761 -34
rect 2551 -114 2761 -94
rect 2475 -942 2481 -166
rect 2515 -942 2521 -166
rect 2475 -954 2521 -942
rect 2633 -166 2679 -154
rect 2633 -942 2639 -166
rect 2673 -942 2679 -166
rect 2633 -1028 2679 -942
rect 2791 -166 2837 14
rect 2867 -34 3077 -14
rect 2867 -94 2887 -34
rect 3057 -94 3077 -34
rect 2867 -114 3077 -94
rect 2791 -942 2797 -166
rect 2831 -942 2837 -166
rect 2791 -954 2837 -942
rect 2949 -166 2995 -154
rect 2949 -942 2955 -166
rect 2989 -942 2995 -166
rect 2949 -1028 2995 -942
rect 3107 -166 3153 14
rect 3183 -34 3283 -14
rect 3183 -94 3203 -34
rect 3263 -94 3283 -34
rect 3183 -114 3283 -94
rect 3107 -942 3113 -166
rect 3147 -942 3153 -166
rect 3107 -954 3153 -942
rect 3265 -166 3471 -154
rect 3265 -942 3271 -166
rect 3305 -184 3471 -166
rect 3305 -924 3411 -184
rect 3451 -924 3471 -184
rect 3305 -942 3471 -924
rect 3265 -1028 3471 -942
rect 261 -1048 3471 -1028
rect 261 -1088 445 -1048
rect 3287 -1088 3471 -1048
rect -554 -1134 168 -1114
rect 261 -1128 3471 -1088
rect 3624 -186 3724 -156
rect 3624 -1104 3644 -186
rect 3684 -1104 3724 -186
rect -554 -1174 -318 -1134
rect 138 -1174 168 -1134
rect -554 -1214 168 -1174
rect 68 -1260 168 -1214
rect 3624 -1260 3724 -1104
rect 68 -1280 3724 -1260
rect 68 -1320 264 -1280
rect 3468 -1320 3724 -1280
rect 68 -1360 3724 -1320
<< via1 >>
rect 599 34 3133 94
rect 127 -96 187 -36
rect 469 -94 529 -34
rect -131 -872 -71 -812
rect 71 -872 131 -812
rect 675 -94 845 -34
rect 991 -94 1161 -34
rect 1307 -94 1477 -34
rect 1623 -94 1793 -34
rect 1939 -94 2109 -34
rect 2255 -94 2425 -34
rect 2571 -94 2741 -34
rect 2887 -94 3057 -34
rect 3203 -94 3263 -34
<< metal2 >>
rect 579 94 3517 114
rect 579 34 599 94
rect 3133 34 3517 94
rect 579 14 3517 34
rect 215 -16 3283 -14
rect 107 -34 3283 -16
rect 107 -36 469 -34
rect 107 -96 127 -36
rect 187 -94 469 -36
rect 529 -94 675 -34
rect 845 -94 991 -34
rect 1161 -94 1307 -34
rect 1477 -94 1623 -34
rect 1793 -94 1939 -34
rect 2109 -94 2255 -34
rect 2425 -94 2571 -34
rect 2741 -94 2887 -34
rect 3057 -94 3203 -34
rect 3263 -94 3283 -34
rect 187 -96 3283 -94
rect 107 -114 3283 -96
rect 107 -116 395 -114
rect -151 -812 -51 -792
rect -151 -872 -131 -812
rect -71 -872 -51 -812
rect -151 -892 -51 -872
rect 51 -812 151 -792
rect 51 -872 71 -812
rect 131 -872 151 -812
rect 51 -892 151 -872
<< labels >>
rlabel metal2 51 -892 151 -792 5 QN
rlabel metal2 -151 -892 -51 -792 5 Q
rlabel metal2 3417 14 3517 114 3 out
rlabel metal1 261 2476 361 2576 1 VDD
rlabel metal1 261 -1128 361 -1028 5 VSS
<< end >>
